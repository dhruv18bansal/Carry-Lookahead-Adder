magic
tech scmos
timestamp 1731689503
<< nwell >>
rect 126 937 167 977
rect 193 937 234 977
rect 248 937 291 977
rect 301 934 331 974
rect 14 -61 44 -21
rect 74 -23 87 -14
rect 74 -63 104 -23
rect 128 -54 158 -14
<< ntransistor >>
rect 139 905 141 915
rect 207 905 209 915
rect 218 905 220 915
rect 262 905 264 915
rect 275 905 277 915
rect 314 909 316 919
rect 27 -86 29 -76
rect 87 -88 89 -78
rect 141 -97 143 -87
<< ptransistor >>
rect 139 943 141 963
rect 151 943 153 963
rect 218 943 220 963
rect 262 943 264 963
rect 314 940 316 960
rect 27 -55 29 -35
rect 87 -57 89 -37
rect 141 -48 143 -28
<< ndiffusion >>
rect 308 915 314 919
rect 133 911 139 915
rect 133 905 134 911
rect 138 905 139 911
rect 141 911 156 915
rect 160 911 161 915
rect 141 905 161 911
rect 200 911 207 915
rect 200 905 201 911
rect 205 905 207 911
rect 209 905 218 915
rect 220 911 223 915
rect 227 911 228 915
rect 220 905 228 911
rect 255 911 262 915
rect 255 905 256 911
rect 260 905 262 911
rect 264 905 275 915
rect 277 911 280 915
rect 284 911 285 915
rect 277 905 285 911
rect 308 909 309 915
rect 313 909 314 915
rect 316 915 318 919
rect 323 915 324 919
rect 316 909 324 915
rect 21 -80 27 -76
rect 21 -86 22 -80
rect 26 -86 27 -80
rect 29 -80 31 -76
rect 36 -80 37 -76
rect 29 -86 37 -80
rect 81 -82 87 -78
rect 81 -88 82 -82
rect 86 -88 87 -82
rect 89 -82 91 -78
rect 96 -82 97 -78
rect 89 -88 97 -82
rect 139 -91 141 -87
rect 135 -97 141 -91
rect 143 -93 151 -87
rect 143 -97 146 -93
<< pdiffusion >>
rect 138 956 139 963
rect 133 943 139 956
rect 141 943 151 963
rect 153 948 161 963
rect 153 943 156 948
rect 160 943 161 948
rect 205 956 218 963
rect 200 943 218 956
rect 220 948 228 963
rect 220 943 223 948
rect 227 943 228 948
rect 260 956 262 963
rect 255 943 262 956
rect 264 948 285 963
rect 264 943 280 948
rect 284 943 285 948
rect 313 953 314 960
rect 308 940 314 953
rect 316 945 324 960
rect 316 940 318 945
rect 323 940 324 945
rect 26 -42 27 -35
rect 21 -55 27 -42
rect 29 -50 37 -35
rect 29 -55 31 -50
rect 36 -55 37 -50
rect 86 -44 87 -37
rect 81 -57 87 -44
rect 89 -52 97 -37
rect 135 -43 141 -28
rect 139 -48 141 -43
rect 143 -33 145 -28
rect 149 -33 151 -28
rect 143 -48 151 -33
rect 89 -57 91 -52
rect 96 -57 97 -52
<< ndcontact >>
rect 134 905 138 911
rect 156 911 160 915
rect 201 905 205 911
rect 223 911 227 915
rect 256 905 260 911
rect 280 911 284 915
rect 309 909 313 915
rect 318 915 323 919
rect 22 -86 26 -80
rect 31 -80 36 -76
rect 82 -88 86 -82
rect 91 -82 96 -78
rect 135 -91 139 -87
rect 146 -97 151 -93
<< pdcontact >>
rect 133 956 138 963
rect 156 943 160 948
rect 200 956 205 963
rect 223 943 227 948
rect 255 956 260 963
rect 280 943 284 948
rect 308 953 313 960
rect 318 940 323 945
rect 21 -42 26 -35
rect 31 -55 36 -50
rect 81 -44 86 -37
rect 135 -48 139 -43
rect 145 -33 149 -28
rect 91 -57 96 -52
<< psubstratepcontact >>
rect 128 891 142 896
rect 148 891 157 896
rect 195 891 209 896
rect 215 891 224 896
rect 250 891 264 896
rect 272 891 281 896
rect 303 895 326 900
rect 16 -100 39 -95
rect 85 -102 99 -97
rect 130 -111 153 -106
<< nsubstratencontact >>
rect 129 970 133 974
rect 137 970 141 974
rect 151 970 155 974
rect 196 970 200 974
rect 204 970 208 974
rect 218 970 222 974
rect 251 970 255 974
rect 259 970 263 974
rect 275 970 279 974
rect 304 967 308 971
rect 312 967 316 971
rect 320 967 324 971
rect 131 -21 135 -17
rect 139 -21 143 -17
rect 147 -21 151 -17
rect 17 -28 21 -24
rect 25 -28 29 -24
rect 33 -28 37 -24
rect 77 -30 81 -26
rect 85 -30 89 -26
rect 93 -30 97 -26
<< polysilicon >>
rect 139 963 141 967
rect 151 963 153 967
rect 218 963 220 967
rect 262 963 264 966
rect 314 960 316 964
rect 139 924 141 943
rect 151 936 153 943
rect 218 936 220 943
rect 152 930 153 936
rect 219 930 220 936
rect 140 919 141 924
rect 151 920 153 930
rect 139 915 141 919
rect 207 915 209 930
rect 218 929 220 930
rect 218 924 220 925
rect 219 919 220 924
rect 262 923 264 943
rect 275 933 277 934
rect 276 927 277 933
rect 314 928 316 940
rect 218 915 220 919
rect 263 917 264 923
rect 262 915 264 917
rect 275 915 277 927
rect 315 923 316 928
rect 314 919 316 923
rect 139 900 141 905
rect 207 902 209 905
rect 218 902 220 905
rect 262 902 264 905
rect 275 902 277 905
rect 314 904 316 909
rect 141 -28 143 -24
rect 27 -35 29 -31
rect 87 -37 89 -33
rect 27 -67 29 -55
rect 141 -57 143 -48
rect 28 -72 29 -67
rect 87 -69 89 -57
rect 141 -62 142 -57
rect 141 -64 143 -62
rect 27 -76 29 -72
rect 88 -74 89 -69
rect 87 -78 89 -74
rect 27 -91 29 -86
rect 141 -79 143 -76
rect 141 -85 142 -79
rect 141 -87 143 -85
rect 87 -93 89 -88
rect 141 -102 143 -97
<< polycontact >>
rect 146 930 152 936
rect 204 930 219 936
rect 134 919 140 924
rect 213 919 219 924
rect 268 927 276 933
rect 254 917 263 923
rect 309 923 315 928
rect 22 -72 28 -67
rect 142 -62 155 -57
rect 82 -74 88 -69
rect 142 -85 150 -79
<< metal1 >>
rect 107 998 245 1004
rect 107 997 182 998
rect 107 936 116 997
rect 126 974 162 977
rect 126 970 129 974
rect 133 970 137 974
rect 141 970 151 974
rect 155 970 162 974
rect 126 969 162 970
rect 133 963 138 969
rect 107 930 146 936
rect 156 924 160 943
rect 177 936 182 997
rect 193 974 229 977
rect 193 970 196 974
rect 200 970 204 974
rect 208 970 218 974
rect 222 970 229 974
rect 193 969 229 970
rect 200 963 205 969
rect 177 930 204 936
rect 128 919 134 924
rect 156 919 213 924
rect 223 923 227 943
rect 237 933 245 998
rect 248 974 286 977
rect 248 970 251 974
rect 255 970 259 974
rect 263 970 275 974
rect 279 970 286 974
rect 248 969 286 970
rect 301 971 331 974
rect 255 963 260 969
rect 301 967 304 971
rect 308 967 312 971
rect 316 967 320 971
rect 324 967 331 971
rect 301 966 331 967
rect 308 960 313 966
rect 237 927 268 933
rect 280 928 284 943
rect 318 928 323 940
rect 280 923 309 928
rect 318 923 335 928
rect 156 915 160 919
rect 223 917 254 923
rect 223 915 227 917
rect 280 915 284 923
rect 318 919 323 923
rect 134 899 138 905
rect 201 899 205 905
rect 256 899 260 905
rect 309 903 313 909
rect 300 900 334 903
rect 125 896 165 899
rect 125 891 128 896
rect 142 891 148 896
rect 157 891 165 896
rect 125 889 165 891
rect 192 896 232 899
rect 192 891 195 896
rect 209 891 215 896
rect 224 891 232 896
rect 192 889 232 891
rect 248 896 289 899
rect 248 891 250 896
rect 264 891 272 896
rect 281 891 289 896
rect 300 895 303 900
rect 326 895 334 900
rect 300 893 334 895
rect 248 889 289 891
rect -3 -67 8 6
rect 65 -2 136 4
rect 14 -24 44 -21
rect 14 -28 17 -24
rect 21 -28 25 -24
rect 29 -28 33 -24
rect 37 -28 44 -24
rect 14 -29 44 -28
rect 21 -35 26 -29
rect -3 -72 22 -67
rect 31 -76 36 -55
rect 65 -69 70 -2
rect 129 -14 136 -2
rect 74 -23 87 -20
rect 128 -17 158 -14
rect 128 -21 131 -17
rect 135 -21 139 -17
rect 143 -21 147 -17
rect 151 -21 158 -17
rect 128 -22 158 -21
rect 74 -26 104 -23
rect 74 -30 77 -26
rect 81 -30 85 -26
rect 89 -30 93 -26
rect 97 -30 104 -26
rect 74 -31 104 -30
rect 145 -28 149 -22
rect 81 -37 86 -31
rect 91 -68 96 -57
rect 135 -68 139 -48
rect 155 -62 166 -57
rect 65 -74 82 -69
rect 91 -72 206 -68
rect 22 -92 26 -86
rect 13 -95 47 -92
rect 13 -100 16 -95
rect 39 -100 47 -95
rect 13 -102 47 -100
rect 65 -112 70 -74
rect 91 -78 96 -72
rect 82 -94 86 -88
rect 135 -87 139 -72
rect 150 -85 174 -79
rect 78 -97 107 -94
rect 78 -100 85 -97
rect 73 -102 85 -100
rect 99 -102 107 -97
rect 73 -104 107 -102
rect 146 -103 151 -97
rect 127 -106 161 -103
rect 127 -111 130 -106
rect 153 -111 161 -106
rect 127 -112 161 -111
rect 65 -113 161 -112
rect 65 -118 134 -113
<< m2contact >>
rect -3 6 8 11
rect 36 -71 41 -66
rect 74 -20 87 -14
rect 166 -62 172 -57
rect 174 -85 187 -79
rect 73 -100 78 -94
<< metal2 >>
rect 8 7 172 11
rect 8 6 87 7
rect 74 -14 87 6
rect 166 -57 172 7
rect 41 -71 64 -66
rect 59 -94 64 -71
rect 59 -100 73 -94
rect 59 -119 67 -100
rect 174 -119 187 -85
rect 59 -128 187 -119
<< labels >>
rlabel metal1 33 -70 33 -70 1 Y
rlabel metal1 42 -100 42 -100 8 gnd
rlabel metal1 33 -23 33 -23 5 vdd
rlabel metal1 201 -71 201 -71 1 out
rlabel metal1 77 -72 77 -72 1 b
rlabel metal1 19 -69 19 -69 1 c
rlabel metal1 160 891 160 891 8 gnd
rlabel metal1 151 975 151 975 5 vdd
rlabel metal1 131 933 133 934 1 clk
rlabel metal1 227 891 227 891 8 gnd
rlabel metal1 218 975 218 975 5 vdd
rlabel metal1 198 933 200 934 1 clk
rlabel metal1 284 891 284 891 8 gnd
rlabel metal1 275 975 275 975 5 vdd
rlabel metal1 329 895 329 895 8 gnd
rlabel metal1 320 972 320 972 5 vdd
rlabel metal1 236 920 240 921 1 1
rlabel metal1 300 926 304 927 1 2
rlabel metal1 129 920 133 922 1 D
rlabel metal1 318 923 321 928 1 Q
<< end >>
