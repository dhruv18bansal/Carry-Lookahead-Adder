magic
tech scmos
timestamp 1731759144
<< nwell >>
rect 1626 -5 1688 22
rect 1722 -10 1749 52
rect 150 -206 212 -179
rect 246 -211 273 -149
rect 721 -196 775 -134
rect 150 -257 212 -230
rect 783 -266 810 -204
rect 1091 -251 1118 -49
rect 1626 -56 1688 -29
rect 1140 -248 1167 -186
rect 1621 -225 1683 -198
rect 1717 -230 1744 -168
rect 1621 -276 1683 -249
rect 163 -355 217 -293
rect 225 -425 252 -363
rect 1081 -866 1135 -804
rect 138 -992 200 -965
rect 234 -997 261 -935
rect 1143 -936 1170 -874
rect 1480 -973 1507 -771
rect 1529 -970 1556 -908
rect 1731 -975 1758 -773
rect 1780 -972 1807 -910
rect 138 -1043 200 -1016
rect 2038 -1035 2100 -1008
rect 2134 -1040 2161 -978
rect 151 -1141 205 -1079
rect 1004 -1111 1058 -1049
rect 1222 -1111 1276 -1049
rect 2038 -1086 2100 -1059
rect -3549 -1226 -3487 -1199
rect -3453 -1231 -3426 -1169
rect -3362 -1247 -3335 -1185
rect -3549 -1277 -3487 -1250
rect -3297 -1344 -3270 -1142
rect -3188 -1216 -3134 -1154
rect 213 -1211 240 -1149
rect 1066 -1181 1093 -1119
rect 1284 -1181 1311 -1119
rect -3248 -1341 -3221 -1279
rect -3126 -1286 -3099 -1224
rect 766 -1403 820 -1341
rect 828 -1473 855 -1411
rect 147 -1652 209 -1625
rect 243 -1657 270 -1595
rect 147 -1703 209 -1676
rect 767 -1686 821 -1624
rect 1003 -1633 1057 -1571
rect 160 -1801 214 -1739
rect 829 -1756 856 -1694
rect 1065 -1703 1092 -1641
rect 1417 -1670 1444 -1468
rect 1466 -1667 1493 -1605
rect 222 -1871 249 -1809
rect 1012 -1844 1066 -1782
rect 763 -1957 817 -1895
rect 1074 -1914 1101 -1852
rect 825 -2027 852 -1965
rect 1428 -1970 1455 -1768
rect 1714 -1823 1741 -1621
rect 2036 -1743 2098 -1716
rect 2132 -1748 2159 -1686
rect 1763 -1820 1790 -1758
rect 2036 -1794 2098 -1767
rect 1477 -1967 1504 -1905
rect 751 -2206 805 -2144
rect 813 -2276 840 -2214
rect 144 -2527 206 -2500
rect 240 -2532 267 -2470
rect 144 -2578 206 -2551
rect 792 -2555 846 -2493
rect 157 -2676 211 -2614
rect 854 -2625 881 -2563
rect 1127 -2607 1181 -2545
rect 1189 -2677 1216 -2615
rect 219 -2746 246 -2684
rect 1457 -2688 1484 -2486
rect 1506 -2685 1533 -2623
rect 2192 -2712 2219 -2510
rect 2241 -2709 2268 -2647
rect 793 -2838 847 -2776
rect 855 -2908 882 -2846
rect 1128 -2890 1182 -2828
rect 1190 -2960 1217 -2898
rect 789 -3109 843 -3047
rect 1464 -3077 1491 -2875
rect 1513 -3074 1540 -3012
rect 851 -3179 878 -3117
rect 1458 -3292 1512 -3230
rect 1756 -3233 1783 -3031
rect 1805 -3230 1832 -3168
rect 777 -3358 831 -3296
rect 1520 -3362 1547 -3300
rect 839 -3428 866 -3366
rect 1118 -3424 1172 -3362
rect 1180 -3494 1207 -3432
rect 794 -3625 848 -3563
rect 856 -3695 883 -3633
rect 782 -3874 836 -3812
rect 844 -3944 871 -3882
<< ntransistor >>
rect 1596 7 1616 9
rect 1699 -5 1701 15
rect 1699 -38 1701 -18
rect 1735 -40 1737 -20
rect 1596 -44 1616 -42
rect 120 -194 140 -192
rect 223 -206 225 -186
rect 223 -239 225 -219
rect 259 -241 261 -221
rect 120 -245 140 -243
rect 753 -262 755 -222
rect 1591 -213 1611 -211
rect 1694 -225 1696 -205
rect 753 -327 755 -287
rect 796 -296 798 -276
rect 1089 -288 1091 -268
rect 1122 -288 1124 -268
rect 1153 -278 1155 -258
rect 1694 -258 1696 -238
rect 1730 -260 1732 -240
rect 1591 -264 1611 -262
rect 195 -421 197 -381
rect 195 -486 197 -446
rect 238 -455 240 -435
rect 1113 -932 1115 -892
rect 108 -980 128 -978
rect 211 -992 213 -972
rect 211 -1025 213 -1005
rect 1113 -997 1115 -957
rect 1156 -966 1158 -946
rect 247 -1027 249 -1007
rect 1478 -1010 1480 -990
rect 1511 -1010 1513 -990
rect 1542 -1000 1544 -980
rect 1729 -1012 1731 -992
rect 1762 -1012 1764 -992
rect 1793 -1002 1795 -982
rect 2008 -1023 2028 -1021
rect 108 -1031 128 -1029
rect 2111 -1035 2113 -1015
rect 2111 -1068 2113 -1048
rect 2147 -1070 2149 -1050
rect 2008 -1074 2028 -1072
rect -3579 -1214 -3559 -1212
rect -3476 -1226 -3474 -1206
rect -3476 -1259 -3474 -1239
rect 183 -1207 185 -1167
rect -3440 -1261 -3438 -1241
rect -3579 -1265 -3559 -1263
rect -3349 -1277 -3347 -1257
rect -3156 -1282 -3154 -1242
rect 1036 -1177 1038 -1137
rect 1254 -1177 1256 -1137
rect 183 -1272 185 -1232
rect 226 -1241 228 -1221
rect 1036 -1242 1038 -1202
rect 1079 -1211 1081 -1191
rect 1254 -1242 1256 -1202
rect 1297 -1211 1299 -1191
rect -3156 -1347 -3154 -1307
rect -3113 -1316 -3111 -1296
rect -3299 -1381 -3297 -1361
rect -3266 -1381 -3264 -1361
rect -3235 -1371 -3233 -1351
rect 798 -1469 800 -1429
rect 798 -1534 800 -1494
rect 841 -1503 843 -1483
rect 117 -1640 137 -1638
rect 220 -1652 222 -1632
rect 220 -1685 222 -1665
rect 256 -1687 258 -1667
rect 117 -1691 137 -1689
rect 799 -1752 801 -1712
rect 1035 -1699 1037 -1659
rect 1415 -1707 1417 -1687
rect 1448 -1707 1450 -1687
rect 1479 -1697 1481 -1677
rect 1035 -1764 1037 -1724
rect 1078 -1733 1080 -1713
rect 192 -1867 194 -1827
rect 799 -1817 801 -1777
rect 842 -1786 844 -1766
rect 192 -1932 194 -1892
rect 235 -1901 237 -1881
rect 1044 -1910 1046 -1870
rect 2006 -1731 2026 -1729
rect 2109 -1743 2111 -1723
rect 2109 -1776 2111 -1756
rect 2145 -1778 2147 -1758
rect 2006 -1782 2026 -1780
rect 1712 -1860 1714 -1840
rect 1745 -1860 1747 -1840
rect 1776 -1850 1778 -1830
rect 795 -2023 797 -1983
rect 1044 -1975 1046 -1935
rect 1087 -1944 1089 -1924
rect 1426 -2007 1428 -1987
rect 1459 -2007 1461 -1987
rect 1490 -1997 1492 -1977
rect 795 -2088 797 -2048
rect 838 -2057 840 -2037
rect 783 -2272 785 -2232
rect 783 -2337 785 -2297
rect 826 -2306 828 -2286
rect 114 -2515 134 -2513
rect 217 -2527 219 -2507
rect 217 -2560 219 -2540
rect 253 -2562 255 -2542
rect 114 -2566 134 -2564
rect 824 -2621 826 -2581
rect 189 -2742 191 -2702
rect 824 -2686 826 -2646
rect 867 -2655 869 -2635
rect 1159 -2673 1161 -2633
rect 1159 -2738 1161 -2698
rect 1202 -2707 1204 -2687
rect 1455 -2725 1457 -2705
rect 1488 -2725 1490 -2705
rect 1519 -2715 1521 -2695
rect 2190 -2749 2192 -2729
rect 2223 -2749 2225 -2729
rect 2254 -2739 2256 -2719
rect 189 -2807 191 -2767
rect 232 -2776 234 -2756
rect 825 -2904 827 -2864
rect 825 -2969 827 -2929
rect 868 -2938 870 -2918
rect 1160 -2956 1162 -2916
rect 1160 -3021 1162 -2981
rect 1203 -2990 1205 -2970
rect 1462 -3114 1464 -3094
rect 1495 -3114 1497 -3094
rect 1526 -3104 1528 -3084
rect 821 -3175 823 -3135
rect 821 -3240 823 -3200
rect 864 -3209 866 -3189
rect 1754 -3270 1756 -3250
rect 1787 -3270 1789 -3250
rect 1818 -3260 1820 -3240
rect 1490 -3358 1492 -3318
rect 809 -3424 811 -3384
rect 809 -3489 811 -3449
rect 852 -3458 854 -3438
rect 1490 -3423 1492 -3383
rect 1533 -3392 1535 -3372
rect 1150 -3490 1152 -3450
rect 1150 -3555 1152 -3515
rect 1193 -3524 1195 -3504
rect 826 -3691 828 -3651
rect 826 -3756 828 -3716
rect 869 -3725 871 -3705
rect 814 -3940 816 -3900
rect 814 -4005 816 -3965
rect 857 -3974 859 -3954
<< ptransistor >>
rect 1634 7 1674 9
rect 1735 -2 1737 38
rect 1634 -44 1674 -42
rect 1104 -143 1106 -63
rect 158 -194 198 -192
rect 259 -203 261 -163
rect 734 -188 736 -148
rect 761 -188 763 -148
rect 158 -245 198 -243
rect 796 -258 798 -218
rect 1104 -243 1106 -163
rect 1153 -240 1155 -200
rect 1629 -213 1669 -211
rect 1730 -222 1732 -182
rect 176 -347 178 -307
rect 203 -347 205 -307
rect 1629 -264 1669 -262
rect 238 -417 240 -377
rect 1094 -858 1096 -818
rect 1121 -858 1123 -818
rect 1493 -865 1495 -785
rect 1744 -867 1746 -787
rect 1156 -928 1158 -888
rect 146 -980 186 -978
rect 247 -989 249 -949
rect 1493 -965 1495 -885
rect 1542 -962 1544 -922
rect 1744 -967 1746 -887
rect 1793 -964 1795 -924
rect 2046 -1023 2086 -1021
rect 146 -1031 186 -1029
rect 2147 -1032 2149 -992
rect 164 -1133 166 -1093
rect 191 -1133 193 -1093
rect 1017 -1103 1019 -1063
rect 1044 -1103 1046 -1063
rect 1235 -1103 1237 -1063
rect 1262 -1103 1264 -1063
rect 2046 -1074 2086 -1072
rect -3541 -1214 -3501 -1212
rect -3440 -1223 -3438 -1183
rect -3349 -1239 -3347 -1199
rect -3284 -1236 -3282 -1156
rect -3175 -1208 -3173 -1168
rect -3148 -1208 -3146 -1168
rect -3541 -1265 -3501 -1263
rect -3284 -1336 -3282 -1256
rect -3235 -1333 -3233 -1293
rect 226 -1203 228 -1163
rect 1079 -1173 1081 -1133
rect -3113 -1278 -3111 -1238
rect 1297 -1173 1299 -1133
rect 779 -1395 781 -1355
rect 806 -1395 808 -1355
rect 841 -1465 843 -1425
rect 1430 -1562 1432 -1482
rect 155 -1640 195 -1638
rect 256 -1649 258 -1609
rect 1016 -1625 1018 -1585
rect 1043 -1625 1045 -1585
rect 780 -1678 782 -1638
rect 807 -1678 809 -1638
rect 155 -1691 195 -1689
rect 173 -1793 175 -1753
rect 200 -1793 202 -1753
rect 842 -1748 844 -1708
rect 1078 -1695 1080 -1655
rect 1430 -1662 1432 -1582
rect 1479 -1659 1481 -1619
rect 1727 -1715 1729 -1635
rect 235 -1863 237 -1823
rect 1025 -1836 1027 -1796
rect 1052 -1836 1054 -1796
rect 776 -1949 778 -1909
rect 803 -1949 805 -1909
rect 1441 -1862 1443 -1782
rect 1727 -1815 1729 -1735
rect 2044 -1731 2084 -1729
rect 2145 -1740 2147 -1700
rect 1776 -1812 1778 -1772
rect 2044 -1782 2084 -1780
rect 1087 -1906 1089 -1866
rect 1441 -1962 1443 -1882
rect 838 -2019 840 -1979
rect 1490 -1959 1492 -1919
rect 764 -2198 766 -2158
rect 791 -2198 793 -2158
rect 826 -2268 828 -2228
rect 152 -2515 192 -2513
rect 253 -2524 255 -2484
rect 805 -2547 807 -2507
rect 832 -2547 834 -2507
rect 152 -2566 192 -2564
rect 170 -2668 172 -2628
rect 197 -2668 199 -2628
rect 867 -2617 869 -2577
rect 1140 -2599 1142 -2559
rect 1167 -2599 1169 -2559
rect 1470 -2580 1472 -2500
rect 1202 -2669 1204 -2629
rect 1470 -2680 1472 -2600
rect 232 -2738 234 -2698
rect 2205 -2604 2207 -2524
rect 1519 -2677 1521 -2637
rect 2205 -2704 2207 -2624
rect 2254 -2701 2256 -2661
rect 806 -2830 808 -2790
rect 833 -2830 835 -2790
rect 868 -2900 870 -2860
rect 1141 -2882 1143 -2842
rect 1168 -2882 1170 -2842
rect 1203 -2952 1205 -2912
rect 1477 -2969 1479 -2889
rect 802 -3101 804 -3061
rect 829 -3101 831 -3061
rect 1477 -3069 1479 -2989
rect 1526 -3066 1528 -3026
rect 1769 -3125 1771 -3045
rect 864 -3171 866 -3131
rect 1769 -3225 1771 -3145
rect 1471 -3284 1473 -3244
rect 1498 -3284 1500 -3244
rect 1818 -3222 1820 -3182
rect 790 -3350 792 -3310
rect 817 -3350 819 -3310
rect 1533 -3354 1535 -3314
rect 852 -3420 854 -3380
rect 1131 -3416 1133 -3376
rect 1158 -3416 1160 -3376
rect 1193 -3486 1195 -3446
rect 807 -3617 809 -3577
rect 834 -3617 836 -3577
rect 869 -3687 871 -3647
rect 795 -3866 797 -3826
rect 822 -3866 824 -3826
rect 857 -3936 859 -3896
<< ndiffusion >>
rect 1596 9 1616 10
rect 1596 6 1616 7
rect 1698 -5 1699 15
rect 1701 -5 1702 15
rect 1596 -42 1616 -41
rect 1698 -38 1699 -18
rect 1701 -38 1702 -18
rect 1734 -40 1735 -20
rect 1737 -40 1738 -20
rect 1596 -45 1616 -44
rect 120 -192 140 -191
rect 120 -195 140 -194
rect 222 -206 223 -186
rect 225 -206 226 -186
rect 120 -243 140 -242
rect 222 -239 223 -219
rect 225 -239 226 -219
rect 258 -241 259 -221
rect 261 -241 262 -221
rect 120 -246 140 -245
rect 752 -262 753 -222
rect 755 -262 756 -222
rect 1591 -211 1611 -210
rect 1591 -214 1611 -213
rect 1693 -225 1694 -205
rect 1696 -225 1697 -205
rect 752 -327 753 -287
rect 755 -327 756 -287
rect 795 -296 796 -276
rect 798 -296 799 -276
rect 1088 -288 1089 -268
rect 1091 -288 1092 -268
rect 1121 -288 1122 -268
rect 1124 -288 1125 -268
rect 1152 -278 1153 -258
rect 1155 -278 1156 -258
rect 1591 -262 1611 -261
rect 1693 -258 1694 -238
rect 1696 -258 1697 -238
rect 1729 -260 1730 -240
rect 1732 -260 1733 -240
rect 1591 -265 1611 -264
rect 194 -421 195 -381
rect 197 -421 198 -381
rect 194 -486 195 -446
rect 197 -486 198 -446
rect 237 -455 238 -435
rect 240 -455 241 -435
rect 1112 -932 1113 -892
rect 1115 -932 1116 -892
rect 108 -978 128 -977
rect 108 -981 128 -980
rect 210 -992 211 -972
rect 213 -992 214 -972
rect 108 -1029 128 -1028
rect 210 -1025 211 -1005
rect 213 -1025 214 -1005
rect 1112 -997 1113 -957
rect 1115 -997 1116 -957
rect 1155 -966 1156 -946
rect 1158 -966 1159 -946
rect 246 -1027 247 -1007
rect 249 -1027 250 -1007
rect 1477 -1010 1478 -990
rect 1480 -1010 1481 -990
rect 1510 -1010 1511 -990
rect 1513 -1010 1514 -990
rect 1541 -1000 1542 -980
rect 1544 -1000 1545 -980
rect 1728 -1012 1729 -992
rect 1731 -1012 1732 -992
rect 1761 -1012 1762 -992
rect 1764 -1012 1765 -992
rect 1792 -1002 1793 -982
rect 1795 -1002 1796 -982
rect 2008 -1021 2028 -1020
rect 2008 -1024 2028 -1023
rect 108 -1032 128 -1031
rect 2110 -1035 2111 -1015
rect 2113 -1035 2114 -1015
rect 2008 -1072 2028 -1071
rect 2110 -1068 2111 -1048
rect 2113 -1068 2114 -1048
rect 2146 -1070 2147 -1050
rect 2149 -1070 2150 -1050
rect 2008 -1075 2028 -1074
rect -3579 -1212 -3559 -1211
rect -3579 -1215 -3559 -1214
rect -3477 -1226 -3476 -1206
rect -3474 -1226 -3473 -1206
rect -3579 -1263 -3559 -1262
rect -3477 -1259 -3476 -1239
rect -3474 -1259 -3473 -1239
rect 182 -1207 183 -1167
rect 185 -1207 186 -1167
rect -3441 -1261 -3440 -1241
rect -3438 -1261 -3437 -1241
rect -3579 -1266 -3559 -1265
rect -3350 -1277 -3349 -1257
rect -3347 -1277 -3346 -1257
rect -3157 -1282 -3156 -1242
rect -3154 -1282 -3153 -1242
rect 1035 -1177 1036 -1137
rect 1038 -1177 1039 -1137
rect 1253 -1177 1254 -1137
rect 1256 -1177 1257 -1137
rect 182 -1272 183 -1232
rect 185 -1272 186 -1232
rect 225 -1241 226 -1221
rect 228 -1241 229 -1221
rect 1035 -1242 1036 -1202
rect 1038 -1242 1039 -1202
rect 1078 -1211 1079 -1191
rect 1081 -1211 1082 -1191
rect 1253 -1242 1254 -1202
rect 1256 -1242 1257 -1202
rect 1296 -1211 1297 -1191
rect 1299 -1211 1300 -1191
rect -3157 -1347 -3156 -1307
rect -3154 -1347 -3153 -1307
rect -3114 -1316 -3113 -1296
rect -3111 -1316 -3110 -1296
rect -3300 -1381 -3299 -1361
rect -3297 -1381 -3296 -1361
rect -3267 -1381 -3266 -1361
rect -3264 -1381 -3263 -1361
rect -3236 -1371 -3235 -1351
rect -3233 -1371 -3232 -1351
rect 797 -1469 798 -1429
rect 800 -1469 801 -1429
rect 797 -1534 798 -1494
rect 800 -1534 801 -1494
rect 840 -1503 841 -1483
rect 843 -1503 844 -1483
rect 117 -1638 137 -1637
rect 117 -1641 137 -1640
rect 219 -1652 220 -1632
rect 222 -1652 223 -1632
rect 117 -1689 137 -1688
rect 219 -1685 220 -1665
rect 222 -1685 223 -1665
rect 255 -1687 256 -1667
rect 258 -1687 259 -1667
rect 117 -1692 137 -1691
rect 798 -1752 799 -1712
rect 801 -1752 802 -1712
rect 1034 -1699 1035 -1659
rect 1037 -1699 1038 -1659
rect 1414 -1707 1415 -1687
rect 1417 -1707 1418 -1687
rect 1447 -1707 1448 -1687
rect 1450 -1707 1451 -1687
rect 1478 -1697 1479 -1677
rect 1481 -1697 1482 -1677
rect 1034 -1764 1035 -1724
rect 1037 -1764 1038 -1724
rect 1077 -1733 1078 -1713
rect 1080 -1733 1081 -1713
rect 191 -1867 192 -1827
rect 194 -1867 195 -1827
rect 798 -1817 799 -1777
rect 801 -1817 802 -1777
rect 841 -1786 842 -1766
rect 844 -1786 845 -1766
rect 191 -1932 192 -1892
rect 194 -1932 195 -1892
rect 234 -1901 235 -1881
rect 237 -1901 238 -1881
rect 1043 -1910 1044 -1870
rect 1046 -1910 1047 -1870
rect 2006 -1729 2026 -1728
rect 2006 -1732 2026 -1731
rect 2108 -1743 2109 -1723
rect 2111 -1743 2112 -1723
rect 2006 -1780 2026 -1779
rect 2108 -1776 2109 -1756
rect 2111 -1776 2112 -1756
rect 2144 -1778 2145 -1758
rect 2147 -1778 2148 -1758
rect 2006 -1783 2026 -1782
rect 1711 -1860 1712 -1840
rect 1714 -1860 1715 -1840
rect 1744 -1860 1745 -1840
rect 1747 -1860 1748 -1840
rect 1775 -1850 1776 -1830
rect 1778 -1850 1779 -1830
rect 794 -2023 795 -1983
rect 797 -2023 798 -1983
rect 1043 -1975 1044 -1935
rect 1046 -1975 1047 -1935
rect 1086 -1944 1087 -1924
rect 1089 -1944 1090 -1924
rect 1425 -2007 1426 -1987
rect 1428 -2007 1429 -1987
rect 1458 -2007 1459 -1987
rect 1461 -2007 1462 -1987
rect 1489 -1997 1490 -1977
rect 1492 -1997 1493 -1977
rect 794 -2088 795 -2048
rect 797 -2088 798 -2048
rect 837 -2057 838 -2037
rect 840 -2057 841 -2037
rect 782 -2272 783 -2232
rect 785 -2272 786 -2232
rect 782 -2337 783 -2297
rect 785 -2337 786 -2297
rect 825 -2306 826 -2286
rect 828 -2306 829 -2286
rect 114 -2513 134 -2512
rect 114 -2516 134 -2515
rect 216 -2527 217 -2507
rect 219 -2527 220 -2507
rect 114 -2564 134 -2563
rect 216 -2560 217 -2540
rect 219 -2560 220 -2540
rect 252 -2562 253 -2542
rect 255 -2562 256 -2542
rect 114 -2567 134 -2566
rect 823 -2621 824 -2581
rect 826 -2621 827 -2581
rect 188 -2742 189 -2702
rect 191 -2742 192 -2702
rect 823 -2686 824 -2646
rect 826 -2686 827 -2646
rect 866 -2655 867 -2635
rect 869 -2655 870 -2635
rect 1158 -2673 1159 -2633
rect 1161 -2673 1162 -2633
rect 1158 -2738 1159 -2698
rect 1161 -2738 1162 -2698
rect 1201 -2707 1202 -2687
rect 1204 -2707 1205 -2687
rect 1454 -2725 1455 -2705
rect 1457 -2725 1458 -2705
rect 1487 -2725 1488 -2705
rect 1490 -2725 1491 -2705
rect 1518 -2715 1519 -2695
rect 1521 -2715 1522 -2695
rect 2189 -2749 2190 -2729
rect 2192 -2749 2193 -2729
rect 2222 -2749 2223 -2729
rect 2225 -2749 2226 -2729
rect 2253 -2739 2254 -2719
rect 2256 -2739 2257 -2719
rect 188 -2807 189 -2767
rect 191 -2807 192 -2767
rect 231 -2776 232 -2756
rect 234 -2776 235 -2756
rect 824 -2904 825 -2864
rect 827 -2904 828 -2864
rect 824 -2969 825 -2929
rect 827 -2969 828 -2929
rect 867 -2938 868 -2918
rect 870 -2938 871 -2918
rect 1159 -2956 1160 -2916
rect 1162 -2956 1163 -2916
rect 1159 -3021 1160 -2981
rect 1162 -3021 1163 -2981
rect 1202 -2990 1203 -2970
rect 1205 -2990 1206 -2970
rect 1461 -3114 1462 -3094
rect 1464 -3114 1465 -3094
rect 1494 -3114 1495 -3094
rect 1497 -3114 1498 -3094
rect 1525 -3104 1526 -3084
rect 1528 -3104 1529 -3084
rect 820 -3175 821 -3135
rect 823 -3175 824 -3135
rect 820 -3240 821 -3200
rect 823 -3240 824 -3200
rect 863 -3209 864 -3189
rect 866 -3209 867 -3189
rect 1753 -3270 1754 -3250
rect 1756 -3270 1757 -3250
rect 1786 -3270 1787 -3250
rect 1789 -3270 1790 -3250
rect 1817 -3260 1818 -3240
rect 1820 -3260 1821 -3240
rect 1489 -3358 1490 -3318
rect 1492 -3358 1493 -3318
rect 808 -3424 809 -3384
rect 811 -3424 812 -3384
rect 808 -3489 809 -3449
rect 811 -3489 812 -3449
rect 851 -3458 852 -3438
rect 854 -3458 855 -3438
rect 1489 -3423 1490 -3383
rect 1492 -3423 1493 -3383
rect 1532 -3392 1533 -3372
rect 1535 -3392 1536 -3372
rect 1149 -3490 1150 -3450
rect 1152 -3490 1153 -3450
rect 1149 -3555 1150 -3515
rect 1152 -3555 1153 -3515
rect 1192 -3524 1193 -3504
rect 1195 -3524 1196 -3504
rect 825 -3691 826 -3651
rect 828 -3691 829 -3651
rect 825 -3756 826 -3716
rect 828 -3756 829 -3716
rect 868 -3725 869 -3705
rect 871 -3725 872 -3705
rect 813 -3940 814 -3900
rect 816 -3940 817 -3900
rect 813 -4005 814 -3965
rect 816 -4005 817 -3965
rect 856 -3974 857 -3954
rect 859 -3974 860 -3954
<< pdiffusion >>
rect 1634 9 1674 10
rect 1634 6 1674 7
rect 1734 -2 1735 38
rect 1737 -2 1738 38
rect 1634 -42 1674 -41
rect 1634 -45 1674 -44
rect 1103 -143 1104 -63
rect 1106 -143 1107 -63
rect 158 -192 198 -191
rect 158 -195 198 -194
rect 258 -203 259 -163
rect 261 -203 262 -163
rect 733 -188 734 -148
rect 736 -188 737 -148
rect 760 -188 761 -148
rect 763 -188 764 -148
rect 158 -243 198 -242
rect 158 -246 198 -245
rect 795 -258 796 -218
rect 798 -258 799 -218
rect 1103 -243 1104 -163
rect 1106 -243 1107 -163
rect 1152 -240 1153 -200
rect 1155 -240 1156 -200
rect 1629 -211 1669 -210
rect 1629 -214 1669 -213
rect 1729 -222 1730 -182
rect 1732 -222 1733 -182
rect 175 -347 176 -307
rect 178 -347 179 -307
rect 202 -347 203 -307
rect 205 -347 206 -307
rect 1629 -262 1669 -261
rect 1629 -265 1669 -264
rect 237 -417 238 -377
rect 240 -417 241 -377
rect 1093 -858 1094 -818
rect 1096 -858 1097 -818
rect 1120 -858 1121 -818
rect 1123 -858 1124 -818
rect 1492 -865 1493 -785
rect 1495 -865 1496 -785
rect 1743 -867 1744 -787
rect 1746 -867 1747 -787
rect 1155 -928 1156 -888
rect 1158 -928 1159 -888
rect 146 -978 186 -977
rect 146 -981 186 -980
rect 246 -989 247 -949
rect 249 -989 250 -949
rect 1492 -965 1493 -885
rect 1495 -965 1496 -885
rect 1541 -962 1542 -922
rect 1544 -962 1545 -922
rect 1743 -967 1744 -887
rect 1746 -967 1747 -887
rect 1792 -964 1793 -924
rect 1795 -964 1796 -924
rect 2046 -1021 2086 -1020
rect 146 -1029 186 -1028
rect 2046 -1024 2086 -1023
rect 146 -1032 186 -1031
rect 2146 -1032 2147 -992
rect 2149 -1032 2150 -992
rect 163 -1133 164 -1093
rect 166 -1133 167 -1093
rect 190 -1133 191 -1093
rect 193 -1133 194 -1093
rect 1016 -1103 1017 -1063
rect 1019 -1103 1020 -1063
rect 1043 -1103 1044 -1063
rect 1046 -1103 1047 -1063
rect 1234 -1103 1235 -1063
rect 1237 -1103 1238 -1063
rect 1261 -1103 1262 -1063
rect 1264 -1103 1265 -1063
rect 2046 -1072 2086 -1071
rect 2046 -1075 2086 -1074
rect -3541 -1212 -3501 -1211
rect -3541 -1215 -3501 -1214
rect -3441 -1223 -3440 -1183
rect -3438 -1223 -3437 -1183
rect -3350 -1239 -3349 -1199
rect -3347 -1239 -3346 -1199
rect -3285 -1236 -3284 -1156
rect -3282 -1236 -3281 -1156
rect -3176 -1208 -3175 -1168
rect -3173 -1208 -3172 -1168
rect -3149 -1208 -3148 -1168
rect -3146 -1208 -3145 -1168
rect -3541 -1263 -3501 -1262
rect -3541 -1266 -3501 -1265
rect -3285 -1336 -3284 -1256
rect -3282 -1336 -3281 -1256
rect -3236 -1333 -3235 -1293
rect -3233 -1333 -3232 -1293
rect 225 -1203 226 -1163
rect 228 -1203 229 -1163
rect 1078 -1173 1079 -1133
rect 1081 -1173 1082 -1133
rect -3114 -1278 -3113 -1238
rect -3111 -1278 -3110 -1238
rect 1296 -1173 1297 -1133
rect 1299 -1173 1300 -1133
rect 778 -1395 779 -1355
rect 781 -1395 782 -1355
rect 805 -1395 806 -1355
rect 808 -1395 809 -1355
rect 840 -1465 841 -1425
rect 843 -1465 844 -1425
rect 1429 -1562 1430 -1482
rect 1432 -1562 1433 -1482
rect 155 -1638 195 -1637
rect 155 -1641 195 -1640
rect 255 -1649 256 -1609
rect 258 -1649 259 -1609
rect 1015 -1625 1016 -1585
rect 1018 -1625 1019 -1585
rect 1042 -1625 1043 -1585
rect 1045 -1625 1046 -1585
rect 779 -1678 780 -1638
rect 782 -1678 783 -1638
rect 806 -1678 807 -1638
rect 809 -1678 810 -1638
rect 155 -1689 195 -1688
rect 155 -1692 195 -1691
rect 172 -1793 173 -1753
rect 175 -1793 176 -1753
rect 199 -1793 200 -1753
rect 202 -1793 203 -1753
rect 841 -1748 842 -1708
rect 844 -1748 845 -1708
rect 1077 -1695 1078 -1655
rect 1080 -1695 1081 -1655
rect 1429 -1662 1430 -1582
rect 1432 -1662 1433 -1582
rect 1478 -1659 1479 -1619
rect 1481 -1659 1482 -1619
rect 1726 -1715 1727 -1635
rect 1729 -1715 1730 -1635
rect 234 -1863 235 -1823
rect 237 -1863 238 -1823
rect 1024 -1836 1025 -1796
rect 1027 -1836 1028 -1796
rect 1051 -1836 1052 -1796
rect 1054 -1836 1055 -1796
rect 775 -1949 776 -1909
rect 778 -1949 779 -1909
rect 802 -1949 803 -1909
rect 805 -1949 806 -1909
rect 1440 -1862 1441 -1782
rect 1443 -1862 1444 -1782
rect 1726 -1815 1727 -1735
rect 1729 -1815 1730 -1735
rect 2044 -1729 2084 -1728
rect 2044 -1732 2084 -1731
rect 2144 -1740 2145 -1700
rect 2147 -1740 2148 -1700
rect 1775 -1812 1776 -1772
rect 1778 -1812 1779 -1772
rect 2044 -1780 2084 -1779
rect 2044 -1783 2084 -1782
rect 1086 -1906 1087 -1866
rect 1089 -1906 1090 -1866
rect 1440 -1962 1441 -1882
rect 1443 -1962 1444 -1882
rect 837 -2019 838 -1979
rect 840 -2019 841 -1979
rect 1489 -1959 1490 -1919
rect 1492 -1959 1493 -1919
rect 763 -2198 764 -2158
rect 766 -2198 767 -2158
rect 790 -2198 791 -2158
rect 793 -2198 794 -2158
rect 825 -2268 826 -2228
rect 828 -2268 829 -2228
rect 152 -2513 192 -2512
rect 152 -2516 192 -2515
rect 252 -2524 253 -2484
rect 255 -2524 256 -2484
rect 804 -2547 805 -2507
rect 807 -2547 808 -2507
rect 831 -2547 832 -2507
rect 834 -2547 835 -2507
rect 152 -2564 192 -2563
rect 152 -2567 192 -2566
rect 169 -2668 170 -2628
rect 172 -2668 173 -2628
rect 196 -2668 197 -2628
rect 199 -2668 200 -2628
rect 866 -2617 867 -2577
rect 869 -2617 870 -2577
rect 1139 -2599 1140 -2559
rect 1142 -2599 1143 -2559
rect 1166 -2599 1167 -2559
rect 1169 -2599 1170 -2559
rect 1469 -2580 1470 -2500
rect 1472 -2580 1473 -2500
rect 1201 -2669 1202 -2629
rect 1204 -2669 1205 -2629
rect 1469 -2680 1470 -2600
rect 1472 -2680 1473 -2600
rect 231 -2738 232 -2698
rect 234 -2738 235 -2698
rect 2204 -2604 2205 -2524
rect 2207 -2604 2208 -2524
rect 1518 -2677 1519 -2637
rect 1521 -2677 1522 -2637
rect 2204 -2704 2205 -2624
rect 2207 -2704 2208 -2624
rect 2253 -2701 2254 -2661
rect 2256 -2701 2257 -2661
rect 805 -2830 806 -2790
rect 808 -2830 809 -2790
rect 832 -2830 833 -2790
rect 835 -2830 836 -2790
rect 867 -2900 868 -2860
rect 870 -2900 871 -2860
rect 1140 -2882 1141 -2842
rect 1143 -2882 1144 -2842
rect 1167 -2882 1168 -2842
rect 1170 -2882 1171 -2842
rect 1202 -2952 1203 -2912
rect 1205 -2952 1206 -2912
rect 1476 -2969 1477 -2889
rect 1479 -2969 1480 -2889
rect 801 -3101 802 -3061
rect 804 -3101 805 -3061
rect 828 -3101 829 -3061
rect 831 -3101 832 -3061
rect 1476 -3069 1477 -2989
rect 1479 -3069 1480 -2989
rect 1525 -3066 1526 -3026
rect 1528 -3066 1529 -3026
rect 1768 -3125 1769 -3045
rect 1771 -3125 1772 -3045
rect 863 -3171 864 -3131
rect 866 -3171 867 -3131
rect 1768 -3225 1769 -3145
rect 1771 -3225 1772 -3145
rect 1470 -3284 1471 -3244
rect 1473 -3284 1474 -3244
rect 1497 -3284 1498 -3244
rect 1500 -3284 1501 -3244
rect 1817 -3222 1818 -3182
rect 1820 -3222 1821 -3182
rect 789 -3350 790 -3310
rect 792 -3350 793 -3310
rect 816 -3350 817 -3310
rect 819 -3350 820 -3310
rect 1532 -3354 1533 -3314
rect 1535 -3354 1536 -3314
rect 851 -3420 852 -3380
rect 854 -3420 855 -3380
rect 1130 -3416 1131 -3376
rect 1133 -3416 1134 -3376
rect 1157 -3416 1158 -3376
rect 1160 -3416 1161 -3376
rect 1192 -3486 1193 -3446
rect 1195 -3486 1196 -3446
rect 806 -3617 807 -3577
rect 809 -3617 810 -3577
rect 833 -3617 834 -3577
rect 836 -3617 837 -3577
rect 868 -3687 869 -3647
rect 871 -3687 872 -3647
rect 794 -3866 795 -3826
rect 797 -3866 798 -3826
rect 821 -3866 822 -3826
rect 824 -3866 825 -3826
rect 856 -3936 857 -3896
rect 859 -3936 860 -3896
<< ndcontact >>
rect 1596 10 1616 14
rect 1596 2 1616 6
rect 1694 -5 1698 15
rect 1702 -5 1706 15
rect 1596 -41 1616 -37
rect 1694 -38 1698 -18
rect 1702 -38 1706 -18
rect 1730 -40 1734 -20
rect 1738 -40 1742 -20
rect 1596 -49 1616 -45
rect 120 -191 140 -187
rect 120 -199 140 -195
rect 218 -206 222 -186
rect 226 -206 230 -186
rect 120 -242 140 -238
rect 218 -239 222 -219
rect 226 -239 230 -219
rect 254 -241 258 -221
rect 262 -241 266 -221
rect 120 -250 140 -246
rect 748 -262 752 -222
rect 756 -262 760 -222
rect 1591 -210 1611 -206
rect 1591 -218 1611 -214
rect 1689 -225 1693 -205
rect 1697 -225 1701 -205
rect 748 -327 752 -287
rect 756 -327 760 -287
rect 791 -296 795 -276
rect 799 -296 803 -276
rect 1084 -288 1088 -268
rect 1092 -288 1096 -268
rect 1117 -288 1121 -268
rect 1125 -288 1129 -268
rect 1148 -278 1152 -258
rect 1156 -278 1160 -258
rect 1591 -261 1611 -257
rect 1689 -258 1693 -238
rect 1697 -258 1701 -238
rect 1725 -260 1729 -240
rect 1733 -260 1737 -240
rect 1591 -269 1611 -265
rect 190 -421 194 -381
rect 198 -421 202 -381
rect 190 -486 194 -446
rect 198 -486 202 -446
rect 233 -455 237 -435
rect 241 -455 245 -435
rect 1108 -932 1112 -892
rect 1116 -932 1120 -892
rect 108 -977 128 -973
rect 108 -985 128 -981
rect 206 -992 210 -972
rect 214 -992 218 -972
rect 108 -1028 128 -1024
rect 206 -1025 210 -1005
rect 214 -1025 218 -1005
rect 1108 -997 1112 -957
rect 1116 -997 1120 -957
rect 1151 -966 1155 -946
rect 1159 -966 1163 -946
rect 242 -1027 246 -1007
rect 250 -1027 254 -1007
rect 1473 -1010 1477 -990
rect 1481 -1010 1485 -990
rect 1506 -1010 1510 -990
rect 1514 -1010 1518 -990
rect 1537 -1000 1541 -980
rect 1545 -1000 1549 -980
rect 1724 -1012 1728 -992
rect 1732 -1012 1736 -992
rect 1757 -1012 1761 -992
rect 1765 -1012 1769 -992
rect 1788 -1002 1792 -982
rect 1796 -1002 1800 -982
rect 2008 -1020 2028 -1016
rect 2008 -1028 2028 -1024
rect 108 -1036 128 -1032
rect 2106 -1035 2110 -1015
rect 2114 -1035 2118 -1015
rect 2008 -1071 2028 -1067
rect 2106 -1068 2110 -1048
rect 2114 -1068 2118 -1048
rect 2142 -1070 2146 -1050
rect 2150 -1070 2154 -1050
rect 2008 -1079 2028 -1075
rect -3579 -1211 -3559 -1207
rect -3579 -1219 -3559 -1215
rect -3481 -1226 -3477 -1206
rect -3473 -1226 -3469 -1206
rect -3579 -1262 -3559 -1258
rect -3481 -1259 -3477 -1239
rect -3473 -1259 -3469 -1239
rect 178 -1207 182 -1167
rect 186 -1207 190 -1167
rect -3445 -1261 -3441 -1241
rect -3437 -1261 -3433 -1241
rect -3579 -1270 -3559 -1266
rect -3354 -1277 -3350 -1257
rect -3346 -1277 -3342 -1257
rect -3161 -1282 -3157 -1242
rect -3153 -1282 -3149 -1242
rect 1031 -1177 1035 -1137
rect 1039 -1177 1043 -1137
rect 1249 -1177 1253 -1137
rect 1257 -1177 1261 -1137
rect 178 -1272 182 -1232
rect 186 -1272 190 -1232
rect 221 -1241 225 -1221
rect 229 -1241 233 -1221
rect 1031 -1242 1035 -1202
rect 1039 -1242 1043 -1202
rect 1074 -1211 1078 -1191
rect 1082 -1211 1086 -1191
rect 1249 -1242 1253 -1202
rect 1257 -1242 1261 -1202
rect 1292 -1211 1296 -1191
rect 1300 -1211 1304 -1191
rect -3161 -1347 -3157 -1307
rect -3153 -1347 -3149 -1307
rect -3118 -1316 -3114 -1296
rect -3110 -1316 -3106 -1296
rect -3304 -1381 -3300 -1361
rect -3296 -1381 -3292 -1361
rect -3271 -1381 -3267 -1361
rect -3263 -1381 -3259 -1361
rect -3240 -1371 -3236 -1351
rect -3232 -1371 -3228 -1351
rect 793 -1469 797 -1429
rect 801 -1469 805 -1429
rect 793 -1534 797 -1494
rect 801 -1534 805 -1494
rect 836 -1503 840 -1483
rect 844 -1503 848 -1483
rect 117 -1637 137 -1633
rect 117 -1645 137 -1641
rect 215 -1652 219 -1632
rect 223 -1652 227 -1632
rect 117 -1688 137 -1684
rect 215 -1685 219 -1665
rect 223 -1685 227 -1665
rect 251 -1687 255 -1667
rect 259 -1687 263 -1667
rect 117 -1696 137 -1692
rect 794 -1752 798 -1712
rect 802 -1752 806 -1712
rect 1030 -1699 1034 -1659
rect 1038 -1699 1042 -1659
rect 1410 -1707 1414 -1687
rect 1418 -1707 1422 -1687
rect 1443 -1707 1447 -1687
rect 1451 -1707 1455 -1687
rect 1474 -1697 1478 -1677
rect 1482 -1697 1486 -1677
rect 1030 -1764 1034 -1724
rect 1038 -1764 1042 -1724
rect 1073 -1733 1077 -1713
rect 1081 -1733 1085 -1713
rect 187 -1867 191 -1827
rect 195 -1867 199 -1827
rect 794 -1817 798 -1777
rect 802 -1817 806 -1777
rect 837 -1786 841 -1766
rect 845 -1786 849 -1766
rect 187 -1932 191 -1892
rect 195 -1932 199 -1892
rect 230 -1901 234 -1881
rect 238 -1901 242 -1881
rect 1039 -1910 1043 -1870
rect 1047 -1910 1051 -1870
rect 2006 -1728 2026 -1724
rect 2006 -1736 2026 -1732
rect 2104 -1743 2108 -1723
rect 2112 -1743 2116 -1723
rect 2006 -1779 2026 -1775
rect 2104 -1776 2108 -1756
rect 2112 -1776 2116 -1756
rect 2140 -1778 2144 -1758
rect 2148 -1778 2152 -1758
rect 2006 -1787 2026 -1783
rect 1707 -1860 1711 -1840
rect 1715 -1860 1719 -1840
rect 1740 -1860 1744 -1840
rect 1748 -1860 1752 -1840
rect 1771 -1850 1775 -1830
rect 1779 -1850 1783 -1830
rect 790 -2023 794 -1983
rect 798 -2023 802 -1983
rect 1039 -1975 1043 -1935
rect 1047 -1975 1051 -1935
rect 1082 -1944 1086 -1924
rect 1090 -1944 1094 -1924
rect 1421 -2007 1425 -1987
rect 1429 -2007 1433 -1987
rect 1454 -2007 1458 -1987
rect 1462 -2007 1466 -1987
rect 1485 -1997 1489 -1977
rect 1493 -1997 1497 -1977
rect 790 -2088 794 -2048
rect 798 -2088 802 -2048
rect 833 -2057 837 -2037
rect 841 -2057 845 -2037
rect 778 -2272 782 -2232
rect 786 -2272 790 -2232
rect 778 -2337 782 -2297
rect 786 -2337 790 -2297
rect 821 -2306 825 -2286
rect 829 -2306 833 -2286
rect 114 -2512 134 -2508
rect 114 -2520 134 -2516
rect 212 -2527 216 -2507
rect 220 -2527 224 -2507
rect 114 -2563 134 -2559
rect 212 -2560 216 -2540
rect 220 -2560 224 -2540
rect 248 -2562 252 -2542
rect 256 -2562 260 -2542
rect 114 -2571 134 -2567
rect 819 -2621 823 -2581
rect 827 -2621 831 -2581
rect 184 -2742 188 -2702
rect 192 -2742 196 -2702
rect 819 -2686 823 -2646
rect 827 -2686 831 -2646
rect 862 -2655 866 -2635
rect 870 -2655 874 -2635
rect 1154 -2673 1158 -2633
rect 1162 -2673 1166 -2633
rect 1154 -2738 1158 -2698
rect 1162 -2738 1166 -2698
rect 1197 -2707 1201 -2687
rect 1205 -2707 1209 -2687
rect 1450 -2725 1454 -2705
rect 1458 -2725 1462 -2705
rect 1483 -2725 1487 -2705
rect 1491 -2725 1495 -2705
rect 1514 -2715 1518 -2695
rect 1522 -2715 1526 -2695
rect 2185 -2749 2189 -2729
rect 2193 -2749 2197 -2729
rect 2218 -2749 2222 -2729
rect 2226 -2749 2230 -2729
rect 2249 -2739 2253 -2719
rect 2257 -2739 2261 -2719
rect 184 -2807 188 -2767
rect 192 -2807 196 -2767
rect 227 -2776 231 -2756
rect 235 -2776 239 -2756
rect 820 -2904 824 -2864
rect 828 -2904 832 -2864
rect 820 -2969 824 -2929
rect 828 -2969 832 -2929
rect 863 -2938 867 -2918
rect 871 -2938 875 -2918
rect 1155 -2956 1159 -2916
rect 1163 -2956 1167 -2916
rect 1155 -3021 1159 -2981
rect 1163 -3021 1167 -2981
rect 1198 -2990 1202 -2970
rect 1206 -2990 1210 -2970
rect 1457 -3114 1461 -3094
rect 1465 -3114 1469 -3094
rect 1490 -3114 1494 -3094
rect 1498 -3114 1502 -3094
rect 1521 -3104 1525 -3084
rect 1529 -3104 1533 -3084
rect 816 -3175 820 -3135
rect 824 -3175 828 -3135
rect 816 -3240 820 -3200
rect 824 -3240 828 -3200
rect 859 -3209 863 -3189
rect 867 -3209 871 -3189
rect 1749 -3270 1753 -3250
rect 1757 -3270 1761 -3250
rect 1782 -3270 1786 -3250
rect 1790 -3270 1794 -3250
rect 1813 -3260 1817 -3240
rect 1821 -3260 1825 -3240
rect 1485 -3358 1489 -3318
rect 1493 -3358 1497 -3318
rect 804 -3424 808 -3384
rect 812 -3424 816 -3384
rect 804 -3489 808 -3449
rect 812 -3489 816 -3449
rect 847 -3458 851 -3438
rect 855 -3458 859 -3438
rect 1485 -3423 1489 -3383
rect 1493 -3423 1497 -3383
rect 1528 -3392 1532 -3372
rect 1536 -3392 1540 -3372
rect 1145 -3490 1149 -3450
rect 1153 -3490 1157 -3450
rect 1145 -3555 1149 -3515
rect 1153 -3555 1157 -3515
rect 1188 -3524 1192 -3504
rect 1196 -3524 1200 -3504
rect 821 -3691 825 -3651
rect 829 -3691 833 -3651
rect 821 -3756 825 -3716
rect 829 -3756 833 -3716
rect 864 -3725 868 -3705
rect 872 -3725 876 -3705
rect 809 -3940 813 -3900
rect 817 -3940 821 -3900
rect 809 -4005 813 -3965
rect 817 -4005 821 -3965
rect 852 -3974 856 -3954
rect 860 -3974 864 -3954
<< pdcontact >>
rect 1634 10 1674 14
rect 1634 2 1674 6
rect 1730 -2 1734 38
rect 1738 -2 1742 38
rect 1634 -41 1674 -37
rect 1634 -49 1674 -45
rect 1099 -143 1103 -63
rect 1107 -143 1111 -63
rect 158 -191 198 -187
rect 158 -199 198 -195
rect 254 -203 258 -163
rect 262 -203 266 -163
rect 729 -188 733 -148
rect 737 -188 741 -148
rect 756 -188 760 -148
rect 764 -188 768 -148
rect 158 -242 198 -238
rect 158 -250 198 -246
rect 791 -258 795 -218
rect 799 -258 803 -218
rect 1099 -243 1103 -163
rect 1107 -243 1111 -163
rect 1148 -240 1152 -200
rect 1156 -240 1160 -200
rect 1629 -210 1669 -206
rect 1629 -218 1669 -214
rect 1725 -222 1729 -182
rect 1733 -222 1737 -182
rect 171 -347 175 -307
rect 179 -347 183 -307
rect 198 -347 202 -307
rect 206 -347 210 -307
rect 1629 -261 1669 -257
rect 1629 -269 1669 -265
rect 233 -417 237 -377
rect 241 -417 245 -377
rect 1089 -858 1093 -818
rect 1097 -858 1101 -818
rect 1116 -858 1120 -818
rect 1124 -858 1128 -818
rect 1488 -865 1492 -785
rect 1496 -865 1500 -785
rect 1739 -867 1743 -787
rect 1747 -867 1751 -787
rect 1151 -928 1155 -888
rect 1159 -928 1163 -888
rect 146 -977 186 -973
rect 146 -985 186 -981
rect 242 -989 246 -949
rect 250 -989 254 -949
rect 146 -1028 186 -1024
rect 1488 -965 1492 -885
rect 1496 -965 1500 -885
rect 1537 -962 1541 -922
rect 1545 -962 1549 -922
rect 1739 -967 1743 -887
rect 1747 -967 1751 -887
rect 1788 -964 1792 -924
rect 1796 -964 1800 -924
rect 2046 -1020 2086 -1016
rect 2046 -1028 2086 -1024
rect 146 -1036 186 -1032
rect 2142 -1032 2146 -992
rect 2150 -1032 2154 -992
rect 159 -1133 163 -1093
rect 167 -1133 171 -1093
rect 186 -1133 190 -1093
rect 194 -1133 198 -1093
rect 1012 -1103 1016 -1063
rect 1020 -1103 1024 -1063
rect 1039 -1103 1043 -1063
rect 1047 -1103 1051 -1063
rect 1230 -1103 1234 -1063
rect 1238 -1103 1242 -1063
rect 1257 -1103 1261 -1063
rect 1265 -1103 1269 -1063
rect 2046 -1071 2086 -1067
rect 2046 -1079 2086 -1075
rect -3541 -1211 -3501 -1207
rect -3541 -1219 -3501 -1215
rect -3445 -1223 -3441 -1183
rect -3437 -1223 -3433 -1183
rect -3541 -1262 -3501 -1258
rect -3354 -1239 -3350 -1199
rect -3346 -1239 -3342 -1199
rect -3289 -1236 -3285 -1156
rect -3281 -1236 -3277 -1156
rect -3180 -1208 -3176 -1168
rect -3172 -1208 -3168 -1168
rect -3153 -1208 -3149 -1168
rect -3145 -1208 -3141 -1168
rect -3541 -1270 -3501 -1266
rect -3289 -1336 -3285 -1256
rect -3281 -1336 -3277 -1256
rect -3240 -1333 -3236 -1293
rect -3232 -1333 -3228 -1293
rect 221 -1203 225 -1163
rect 229 -1203 233 -1163
rect 1074 -1173 1078 -1133
rect 1082 -1173 1086 -1133
rect -3118 -1278 -3114 -1238
rect -3110 -1278 -3106 -1238
rect 1292 -1173 1296 -1133
rect 1300 -1173 1304 -1133
rect 774 -1395 778 -1355
rect 782 -1395 786 -1355
rect 801 -1395 805 -1355
rect 809 -1395 813 -1355
rect 836 -1465 840 -1425
rect 844 -1465 848 -1425
rect 1425 -1562 1429 -1482
rect 1433 -1562 1437 -1482
rect 155 -1637 195 -1633
rect 155 -1645 195 -1641
rect 251 -1649 255 -1609
rect 259 -1649 263 -1609
rect 1011 -1625 1015 -1585
rect 1019 -1625 1023 -1585
rect 1038 -1625 1042 -1585
rect 1046 -1625 1050 -1585
rect 155 -1688 195 -1684
rect 775 -1678 779 -1638
rect 783 -1678 787 -1638
rect 802 -1678 806 -1638
rect 810 -1678 814 -1638
rect 155 -1696 195 -1692
rect 168 -1793 172 -1753
rect 176 -1793 180 -1753
rect 195 -1793 199 -1753
rect 203 -1793 207 -1753
rect 837 -1748 841 -1708
rect 845 -1748 849 -1708
rect 1073 -1695 1077 -1655
rect 1081 -1695 1085 -1655
rect 1425 -1662 1429 -1582
rect 1433 -1662 1437 -1582
rect 1474 -1659 1478 -1619
rect 1482 -1659 1486 -1619
rect 1722 -1715 1726 -1635
rect 1730 -1715 1734 -1635
rect 230 -1863 234 -1823
rect 238 -1863 242 -1823
rect 1020 -1836 1024 -1796
rect 1028 -1836 1032 -1796
rect 1047 -1836 1051 -1796
rect 1055 -1836 1059 -1796
rect 771 -1949 775 -1909
rect 779 -1949 783 -1909
rect 798 -1949 802 -1909
rect 806 -1949 810 -1909
rect 1436 -1862 1440 -1782
rect 1444 -1862 1448 -1782
rect 1722 -1815 1726 -1735
rect 1730 -1815 1734 -1735
rect 2044 -1728 2084 -1724
rect 2044 -1736 2084 -1732
rect 2140 -1740 2144 -1700
rect 2148 -1740 2152 -1700
rect 1771 -1812 1775 -1772
rect 1779 -1812 1783 -1772
rect 2044 -1779 2084 -1775
rect 2044 -1787 2084 -1783
rect 1082 -1906 1086 -1866
rect 1090 -1906 1094 -1866
rect 1436 -1962 1440 -1882
rect 1444 -1962 1448 -1882
rect 833 -2019 837 -1979
rect 841 -2019 845 -1979
rect 1485 -1959 1489 -1919
rect 1493 -1959 1497 -1919
rect 759 -2198 763 -2158
rect 767 -2198 771 -2158
rect 786 -2198 790 -2158
rect 794 -2198 798 -2158
rect 821 -2268 825 -2228
rect 829 -2268 833 -2228
rect 152 -2512 192 -2508
rect 152 -2520 192 -2516
rect 248 -2524 252 -2484
rect 256 -2524 260 -2484
rect 152 -2563 192 -2559
rect 800 -2547 804 -2507
rect 808 -2547 812 -2507
rect 827 -2547 831 -2507
rect 835 -2547 839 -2507
rect 152 -2571 192 -2567
rect 165 -2668 169 -2628
rect 173 -2668 177 -2628
rect 192 -2668 196 -2628
rect 200 -2668 204 -2628
rect 862 -2617 866 -2577
rect 870 -2617 874 -2577
rect 1135 -2599 1139 -2559
rect 1143 -2599 1147 -2559
rect 1162 -2599 1166 -2559
rect 1170 -2599 1174 -2559
rect 1465 -2580 1469 -2500
rect 1473 -2580 1477 -2500
rect 1197 -2669 1201 -2629
rect 1205 -2669 1209 -2629
rect 1465 -2680 1469 -2600
rect 1473 -2680 1477 -2600
rect 227 -2738 231 -2698
rect 235 -2738 239 -2698
rect 2200 -2604 2204 -2524
rect 2208 -2604 2212 -2524
rect 1514 -2677 1518 -2637
rect 1522 -2677 1526 -2637
rect 2200 -2704 2204 -2624
rect 2208 -2704 2212 -2624
rect 2249 -2701 2253 -2661
rect 2257 -2701 2261 -2661
rect 801 -2830 805 -2790
rect 809 -2830 813 -2790
rect 828 -2830 832 -2790
rect 836 -2830 840 -2790
rect 863 -2900 867 -2860
rect 871 -2900 875 -2860
rect 1136 -2882 1140 -2842
rect 1144 -2882 1148 -2842
rect 1163 -2882 1167 -2842
rect 1171 -2882 1175 -2842
rect 1198 -2952 1202 -2912
rect 1206 -2952 1210 -2912
rect 1472 -2969 1476 -2889
rect 1480 -2969 1484 -2889
rect 797 -3101 801 -3061
rect 805 -3101 809 -3061
rect 824 -3101 828 -3061
rect 832 -3101 836 -3061
rect 1472 -3069 1476 -2989
rect 1480 -3069 1484 -2989
rect 1521 -3066 1525 -3026
rect 1529 -3066 1533 -3026
rect 1764 -3125 1768 -3045
rect 1772 -3125 1776 -3045
rect 859 -3171 863 -3131
rect 867 -3171 871 -3131
rect 1764 -3225 1768 -3145
rect 1772 -3225 1776 -3145
rect 1466 -3284 1470 -3244
rect 1474 -3284 1478 -3244
rect 1493 -3284 1497 -3244
rect 1501 -3284 1505 -3244
rect 1813 -3222 1817 -3182
rect 1821 -3222 1825 -3182
rect 785 -3350 789 -3310
rect 793 -3350 797 -3310
rect 812 -3350 816 -3310
rect 820 -3350 824 -3310
rect 1528 -3354 1532 -3314
rect 1536 -3354 1540 -3314
rect 847 -3420 851 -3380
rect 855 -3420 859 -3380
rect 1126 -3416 1130 -3376
rect 1134 -3416 1138 -3376
rect 1153 -3416 1157 -3376
rect 1161 -3416 1165 -3376
rect 1188 -3486 1192 -3446
rect 1196 -3486 1200 -3446
rect 802 -3617 806 -3577
rect 810 -3617 814 -3577
rect 829 -3617 833 -3577
rect 837 -3617 841 -3577
rect 864 -3687 868 -3647
rect 872 -3687 876 -3647
rect 790 -3866 794 -3826
rect 798 -3866 802 -3826
rect 817 -3866 821 -3826
rect 825 -3866 829 -3826
rect 852 -3936 856 -3896
rect 860 -3936 864 -3896
<< psubstratepcontact >>
rect 1585 17 1589 21
rect 1585 -4 1589 0
rect 1585 -34 1589 -30
rect 1585 -55 1589 -51
rect 1723 -51 1727 -47
rect 1744 -51 1748 -47
rect 109 -184 113 -180
rect 109 -205 113 -201
rect 109 -235 113 -231
rect 109 -256 113 -252
rect 247 -252 251 -248
rect 268 -252 272 -248
rect 1580 -203 1584 -199
rect 1580 -224 1584 -220
rect 1580 -254 1584 -250
rect 1580 -275 1584 -271
rect 1718 -271 1722 -267
rect 1739 -271 1743 -267
rect 1141 -289 1145 -285
rect 1162 -289 1166 -285
rect 1077 -299 1081 -295
rect 1098 -299 1102 -295
rect 1110 -299 1114 -295
rect 1131 -299 1135 -295
rect 784 -307 788 -303
rect 805 -307 809 -303
rect 741 -338 745 -334
rect 762 -338 766 -334
rect 226 -466 230 -462
rect 247 -466 251 -462
rect 183 -497 187 -493
rect 204 -497 208 -493
rect 97 -970 101 -966
rect 97 -991 101 -987
rect 97 -1021 101 -1017
rect 1144 -977 1148 -973
rect 1165 -977 1169 -973
rect 1101 -1008 1105 -1004
rect 1122 -1008 1126 -1004
rect 1530 -1011 1534 -1007
rect 1551 -1011 1555 -1007
rect 1781 -1013 1785 -1009
rect 1802 -1013 1806 -1009
rect 1997 -1013 2001 -1009
rect 1466 -1021 1470 -1017
rect 1487 -1021 1491 -1017
rect 1499 -1021 1503 -1017
rect 1520 -1021 1524 -1017
rect 1717 -1023 1721 -1019
rect 1738 -1023 1742 -1019
rect 1750 -1023 1754 -1019
rect 1771 -1023 1775 -1019
rect 1997 -1034 2001 -1030
rect 97 -1042 101 -1038
rect 235 -1038 239 -1034
rect 256 -1038 260 -1034
rect 1997 -1064 2001 -1060
rect 1997 -1085 2001 -1081
rect 2135 -1081 2139 -1077
rect 2156 -1081 2160 -1077
rect -3590 -1204 -3586 -1200
rect -3590 -1225 -3586 -1221
rect -3590 -1255 -3586 -1251
rect -3590 -1276 -3586 -1272
rect -3452 -1272 -3448 -1268
rect -3431 -1272 -3427 -1268
rect -3361 -1288 -3357 -1284
rect -3340 -1288 -3336 -1284
rect 1067 -1222 1071 -1218
rect 1088 -1222 1092 -1218
rect 1285 -1222 1289 -1218
rect 1306 -1222 1310 -1218
rect 214 -1252 218 -1248
rect 235 -1252 239 -1248
rect 1024 -1253 1028 -1249
rect 1045 -1253 1049 -1249
rect 1242 -1253 1246 -1249
rect 1263 -1253 1267 -1249
rect 171 -1283 175 -1279
rect 192 -1283 196 -1279
rect -3125 -1327 -3121 -1323
rect -3104 -1327 -3100 -1323
rect -3168 -1358 -3164 -1354
rect -3147 -1358 -3143 -1354
rect -3247 -1382 -3243 -1378
rect -3226 -1382 -3222 -1378
rect -3311 -1392 -3307 -1388
rect -3290 -1392 -3286 -1388
rect -3278 -1392 -3274 -1388
rect -3257 -1392 -3253 -1388
rect 829 -1514 833 -1510
rect 850 -1514 854 -1510
rect 786 -1545 790 -1541
rect 807 -1545 811 -1541
rect 106 -1630 110 -1626
rect 106 -1651 110 -1647
rect 106 -1681 110 -1677
rect 106 -1702 110 -1698
rect 244 -1698 248 -1694
rect 265 -1698 269 -1694
rect 1467 -1708 1471 -1704
rect 1488 -1708 1492 -1704
rect 1403 -1718 1407 -1714
rect 1424 -1718 1428 -1714
rect 1436 -1718 1440 -1714
rect 1457 -1718 1461 -1714
rect 1995 -1721 1999 -1717
rect 1066 -1744 1070 -1740
rect 1087 -1744 1091 -1740
rect 1023 -1775 1027 -1771
rect 1044 -1775 1048 -1771
rect 830 -1797 834 -1793
rect 851 -1797 855 -1793
rect 787 -1828 791 -1824
rect 808 -1828 812 -1824
rect 223 -1912 227 -1908
rect 244 -1912 248 -1908
rect 180 -1943 184 -1939
rect 201 -1943 205 -1939
rect 1995 -1742 1999 -1738
rect 1995 -1772 1999 -1768
rect 1995 -1793 1999 -1789
rect 2133 -1789 2137 -1785
rect 2154 -1789 2158 -1785
rect 1764 -1861 1768 -1857
rect 1785 -1861 1789 -1857
rect 1075 -1955 1079 -1951
rect 1096 -1955 1100 -1951
rect 1032 -1986 1036 -1982
rect 1053 -1986 1057 -1982
rect 1700 -1871 1704 -1867
rect 1721 -1871 1725 -1867
rect 1733 -1871 1737 -1867
rect 1754 -1871 1758 -1867
rect 1478 -2008 1482 -2004
rect 1499 -2008 1503 -2004
rect 1414 -2018 1418 -2014
rect 1435 -2018 1439 -2014
rect 1447 -2018 1451 -2014
rect 1468 -2018 1472 -2014
rect 826 -2068 830 -2064
rect 847 -2068 851 -2064
rect 783 -2099 787 -2095
rect 804 -2099 808 -2095
rect 814 -2317 818 -2313
rect 835 -2317 839 -2313
rect 771 -2348 775 -2344
rect 792 -2348 796 -2344
rect 103 -2505 107 -2501
rect 103 -2526 107 -2522
rect 103 -2556 107 -2552
rect 103 -2577 107 -2573
rect 241 -2573 245 -2569
rect 262 -2573 266 -2569
rect 855 -2666 859 -2662
rect 876 -2666 880 -2662
rect 812 -2697 816 -2693
rect 833 -2697 837 -2693
rect 1190 -2718 1194 -2714
rect 1211 -2718 1215 -2714
rect 1507 -2726 1511 -2722
rect 1528 -2726 1532 -2722
rect 1443 -2736 1447 -2732
rect 1464 -2736 1468 -2732
rect 1476 -2736 1480 -2732
rect 1497 -2736 1501 -2732
rect 1147 -2749 1151 -2745
rect 1168 -2749 1172 -2745
rect 2242 -2750 2246 -2746
rect 2263 -2750 2267 -2746
rect 2178 -2760 2182 -2756
rect 2199 -2760 2203 -2756
rect 2211 -2760 2215 -2756
rect 2232 -2760 2236 -2756
rect 220 -2787 224 -2783
rect 241 -2787 245 -2783
rect 177 -2818 181 -2814
rect 198 -2818 202 -2814
rect 856 -2949 860 -2945
rect 877 -2949 881 -2945
rect 813 -2980 817 -2976
rect 834 -2980 838 -2976
rect 1191 -3001 1195 -2997
rect 1212 -3001 1216 -2997
rect 1148 -3032 1152 -3028
rect 1169 -3032 1173 -3028
rect 1514 -3115 1518 -3111
rect 1535 -3115 1539 -3111
rect 1450 -3125 1454 -3121
rect 1471 -3125 1475 -3121
rect 1483 -3125 1487 -3121
rect 1504 -3125 1508 -3121
rect 852 -3220 856 -3216
rect 873 -3220 877 -3216
rect 809 -3251 813 -3247
rect 830 -3251 834 -3247
rect 1806 -3271 1810 -3267
rect 1827 -3271 1831 -3267
rect 1742 -3281 1746 -3277
rect 1763 -3281 1767 -3277
rect 1775 -3281 1779 -3277
rect 1796 -3281 1800 -3277
rect 1521 -3403 1525 -3399
rect 1542 -3403 1546 -3399
rect 840 -3469 844 -3465
rect 861 -3469 865 -3465
rect 797 -3500 801 -3496
rect 818 -3500 822 -3496
rect 1478 -3434 1482 -3430
rect 1499 -3434 1503 -3430
rect 1181 -3535 1185 -3531
rect 1202 -3535 1206 -3531
rect 1138 -3566 1142 -3562
rect 1159 -3566 1163 -3562
rect 857 -3736 861 -3732
rect 878 -3736 882 -3732
rect 814 -3767 818 -3763
rect 835 -3767 839 -3763
rect 845 -3985 849 -3981
rect 866 -3985 870 -3981
rect 802 -4016 806 -4012
rect 823 -4016 827 -4012
<< nsubstratencontact >>
rect 1725 45 1729 49
rect 1742 45 1746 49
rect 1681 15 1685 19
rect 1681 -2 1685 2
rect 1681 -36 1685 -32
rect 1094 -56 1098 -52
rect 1111 -56 1115 -52
rect 1681 -53 1685 -49
rect 724 -141 728 -137
rect 741 -141 745 -137
rect 751 -141 755 -137
rect 768 -141 772 -137
rect 249 -156 253 -152
rect 266 -156 270 -152
rect 205 -186 209 -182
rect 205 -203 209 -199
rect 205 -237 209 -233
rect 205 -254 209 -250
rect 786 -211 790 -207
rect 803 -211 807 -207
rect 1720 -175 1724 -171
rect 1737 -175 1741 -171
rect 1143 -193 1147 -189
rect 1160 -193 1164 -189
rect 1676 -205 1680 -201
rect 1676 -222 1680 -218
rect 1676 -256 1680 -252
rect 166 -300 170 -296
rect 183 -300 187 -296
rect 193 -300 197 -296
rect 210 -300 214 -296
rect 1676 -273 1680 -269
rect 228 -370 232 -366
rect 245 -370 249 -366
rect 1483 -778 1487 -774
rect 1500 -778 1504 -774
rect 1734 -780 1738 -776
rect 1751 -780 1755 -776
rect 1084 -811 1088 -807
rect 1101 -811 1105 -807
rect 1111 -811 1115 -807
rect 1128 -811 1132 -807
rect 237 -942 241 -938
rect 254 -942 258 -938
rect 1146 -881 1150 -877
rect 1163 -881 1167 -877
rect 193 -972 197 -968
rect 193 -989 197 -985
rect 193 -1023 197 -1019
rect 1532 -915 1536 -911
rect 1549 -915 1553 -911
rect 1783 -917 1787 -913
rect 1800 -917 1804 -913
rect 2137 -985 2141 -981
rect 2154 -985 2158 -981
rect 2093 -1015 2097 -1011
rect 2093 -1032 2097 -1028
rect 193 -1040 197 -1036
rect 1007 -1056 1011 -1052
rect 1024 -1056 1028 -1052
rect 1034 -1056 1038 -1052
rect 1051 -1056 1055 -1052
rect 1225 -1056 1229 -1052
rect 1242 -1056 1246 -1052
rect 1252 -1056 1256 -1052
rect 1269 -1056 1273 -1052
rect 154 -1086 158 -1082
rect 171 -1086 175 -1082
rect 181 -1086 185 -1082
rect 198 -1086 202 -1082
rect 2093 -1066 2097 -1062
rect 2093 -1083 2097 -1079
rect -3294 -1149 -3290 -1145
rect -3277 -1149 -3273 -1145
rect -3450 -1176 -3446 -1172
rect -3433 -1176 -3429 -1172
rect -3494 -1206 -3490 -1202
rect -3494 -1223 -3490 -1219
rect -3359 -1192 -3355 -1188
rect -3342 -1192 -3338 -1188
rect -3494 -1257 -3490 -1253
rect -3185 -1161 -3181 -1157
rect -3168 -1161 -3164 -1157
rect -3158 -1161 -3154 -1157
rect -3141 -1161 -3137 -1157
rect -3494 -1274 -3490 -1270
rect -3245 -1286 -3241 -1282
rect -3228 -1286 -3224 -1282
rect 216 -1156 220 -1152
rect 233 -1156 237 -1152
rect 1069 -1126 1073 -1122
rect 1086 -1126 1090 -1122
rect -3123 -1231 -3119 -1227
rect -3106 -1231 -3102 -1227
rect 1287 -1126 1291 -1122
rect 1304 -1126 1308 -1122
rect 769 -1348 773 -1344
rect 786 -1348 790 -1344
rect 796 -1348 800 -1344
rect 813 -1348 817 -1344
rect 831 -1418 835 -1414
rect 848 -1418 852 -1414
rect 1420 -1475 1424 -1471
rect 1437 -1475 1441 -1471
rect 1006 -1578 1010 -1574
rect 1023 -1578 1027 -1574
rect 1033 -1578 1037 -1574
rect 1050 -1578 1054 -1574
rect 246 -1602 250 -1598
rect 263 -1602 267 -1598
rect 202 -1632 206 -1628
rect 202 -1649 206 -1645
rect 770 -1631 774 -1627
rect 787 -1631 791 -1627
rect 797 -1631 801 -1627
rect 814 -1631 818 -1627
rect 202 -1683 206 -1679
rect 202 -1700 206 -1696
rect 163 -1746 167 -1742
rect 180 -1746 184 -1742
rect 190 -1746 194 -1742
rect 207 -1746 211 -1742
rect 832 -1701 836 -1697
rect 849 -1701 853 -1697
rect 1068 -1648 1072 -1644
rect 1085 -1648 1089 -1644
rect 1469 -1612 1473 -1608
rect 1486 -1612 1490 -1608
rect 1717 -1628 1721 -1624
rect 1734 -1628 1738 -1624
rect 2135 -1693 2139 -1689
rect 2152 -1693 2156 -1689
rect 2091 -1723 2095 -1719
rect 225 -1816 229 -1812
rect 242 -1816 246 -1812
rect 1431 -1775 1435 -1771
rect 1448 -1775 1452 -1771
rect 1015 -1789 1019 -1785
rect 1032 -1789 1036 -1785
rect 1042 -1789 1046 -1785
rect 1059 -1789 1063 -1785
rect 766 -1902 770 -1898
rect 783 -1902 787 -1898
rect 793 -1902 797 -1898
rect 810 -1902 814 -1898
rect 1077 -1859 1081 -1855
rect 1094 -1859 1098 -1855
rect 2091 -1740 2095 -1736
rect 1766 -1765 1770 -1761
rect 1783 -1765 1787 -1761
rect 2091 -1774 2095 -1770
rect 2091 -1791 2095 -1787
rect 828 -1972 832 -1968
rect 845 -1972 849 -1968
rect 1480 -1912 1484 -1908
rect 1497 -1912 1501 -1908
rect 754 -2151 758 -2147
rect 771 -2151 775 -2147
rect 781 -2151 785 -2147
rect 798 -2151 802 -2147
rect 816 -2221 820 -2217
rect 833 -2221 837 -2217
rect 243 -2477 247 -2473
rect 260 -2477 264 -2473
rect 199 -2507 203 -2503
rect 199 -2524 203 -2520
rect 1460 -2493 1464 -2489
rect 1477 -2493 1481 -2489
rect 795 -2500 799 -2496
rect 812 -2500 816 -2496
rect 822 -2500 826 -2496
rect 839 -2500 843 -2496
rect 199 -2558 203 -2554
rect 199 -2575 203 -2571
rect 1130 -2552 1134 -2548
rect 1147 -2552 1151 -2548
rect 1157 -2552 1161 -2548
rect 1174 -2552 1178 -2548
rect 160 -2621 164 -2617
rect 177 -2621 181 -2617
rect 187 -2621 191 -2617
rect 204 -2621 208 -2617
rect 857 -2570 861 -2566
rect 874 -2570 878 -2566
rect 2195 -2517 2199 -2513
rect 2212 -2517 2216 -2513
rect 222 -2691 226 -2687
rect 239 -2691 243 -2687
rect 1192 -2622 1196 -2618
rect 1209 -2622 1213 -2618
rect 1509 -2630 1513 -2626
rect 1526 -2630 1530 -2626
rect 2244 -2654 2248 -2650
rect 2261 -2654 2265 -2650
rect 796 -2783 800 -2779
rect 813 -2783 817 -2779
rect 823 -2783 827 -2779
rect 840 -2783 844 -2779
rect 1131 -2835 1135 -2831
rect 1148 -2835 1152 -2831
rect 1158 -2835 1162 -2831
rect 1175 -2835 1179 -2831
rect 858 -2853 862 -2849
rect 875 -2853 879 -2849
rect 1467 -2882 1471 -2878
rect 1484 -2882 1488 -2878
rect 1193 -2905 1197 -2901
rect 1210 -2905 1214 -2901
rect 792 -3054 796 -3050
rect 809 -3054 813 -3050
rect 819 -3054 823 -3050
rect 836 -3054 840 -3050
rect 1516 -3019 1520 -3015
rect 1533 -3019 1537 -3015
rect 1759 -3038 1763 -3034
rect 1776 -3038 1780 -3034
rect 854 -3124 858 -3120
rect 871 -3124 875 -3120
rect 1461 -3237 1465 -3233
rect 1478 -3237 1482 -3233
rect 1488 -3237 1492 -3233
rect 1505 -3237 1509 -3233
rect 1808 -3175 1812 -3171
rect 1825 -3175 1829 -3171
rect 780 -3303 784 -3299
rect 797 -3303 801 -3299
rect 807 -3303 811 -3299
rect 824 -3303 828 -3299
rect 1121 -3369 1125 -3365
rect 1138 -3369 1142 -3365
rect 1148 -3369 1152 -3365
rect 1165 -3369 1169 -3365
rect 842 -3373 846 -3369
rect 859 -3373 863 -3369
rect 1523 -3307 1527 -3303
rect 1540 -3307 1544 -3303
rect 1183 -3439 1187 -3435
rect 1200 -3439 1204 -3435
rect 797 -3570 801 -3566
rect 814 -3570 818 -3566
rect 824 -3570 828 -3566
rect 841 -3570 845 -3566
rect 859 -3640 863 -3636
rect 876 -3640 880 -3636
rect 785 -3819 789 -3815
rect 802 -3819 806 -3815
rect 812 -3819 816 -3815
rect 829 -3819 833 -3815
rect 847 -3889 851 -3885
rect 864 -3889 868 -3885
<< polysilicon >>
rect 1619 37 1701 39
rect 1735 38 1737 41
rect 1699 15 1701 37
rect 1593 7 1596 9
rect 1616 7 1634 9
rect 1674 7 1677 9
rect 1699 -8 1701 -5
rect 1619 -15 1701 -13
rect 1699 -18 1701 -15
rect 1735 -20 1737 -2
rect 1699 -41 1701 -38
rect 1593 -44 1596 -42
rect 1616 -44 1634 -42
rect 1674 -44 1677 -42
rect 1735 -43 1737 -40
rect 1104 -63 1106 -60
rect 734 -148 736 -145
rect 761 -148 763 -145
rect 143 -164 225 -162
rect 259 -163 261 -160
rect 223 -186 225 -164
rect 117 -194 120 -192
rect 140 -194 158 -192
rect 198 -194 201 -192
rect 1104 -149 1106 -143
rect 1104 -151 1124 -149
rect 1104 -163 1106 -160
rect 223 -209 225 -206
rect 143 -216 225 -214
rect 223 -219 225 -216
rect 259 -221 261 -203
rect 734 -216 736 -188
rect 761 -200 763 -188
rect 761 -202 771 -200
rect 734 -218 755 -216
rect 223 -242 225 -239
rect 753 -222 755 -218
rect 117 -245 120 -243
rect 140 -245 158 -243
rect 198 -245 201 -243
rect 259 -244 261 -241
rect 753 -266 755 -262
rect 769 -279 771 -202
rect 796 -218 798 -215
rect 1104 -249 1106 -243
rect 1089 -251 1106 -249
rect 796 -276 798 -258
rect 1089 -268 1091 -251
rect 1122 -268 1124 -151
rect 1614 -183 1696 -181
rect 1730 -182 1732 -179
rect 1153 -200 1155 -197
rect 1694 -205 1696 -183
rect 1588 -213 1591 -211
rect 1611 -213 1629 -211
rect 1669 -213 1672 -211
rect 1694 -228 1696 -225
rect 1614 -235 1696 -233
rect 1694 -238 1696 -235
rect 1153 -258 1155 -240
rect 753 -281 771 -279
rect 753 -287 755 -281
rect 176 -307 178 -304
rect 203 -307 205 -304
rect 1730 -240 1732 -222
rect 1694 -261 1696 -258
rect 1588 -264 1591 -262
rect 1611 -264 1629 -262
rect 1669 -264 1672 -262
rect 1730 -263 1732 -260
rect 1153 -281 1155 -278
rect 1089 -291 1091 -288
rect 1122 -291 1124 -288
rect 796 -299 798 -296
rect 753 -330 755 -327
rect 176 -375 178 -347
rect 203 -359 205 -347
rect 203 -361 213 -359
rect 176 -377 197 -375
rect 195 -381 197 -377
rect 195 -425 197 -421
rect 211 -438 213 -361
rect 238 -377 240 -374
rect 238 -435 240 -417
rect 195 -440 213 -438
rect 195 -446 197 -440
rect 238 -458 240 -455
rect 195 -489 197 -486
rect 1493 -785 1495 -782
rect 1094 -818 1096 -815
rect 1121 -818 1123 -815
rect 1094 -886 1096 -858
rect 1121 -870 1123 -858
rect 1744 -787 1746 -784
rect 1121 -872 1131 -870
rect 1094 -888 1115 -886
rect 1113 -892 1115 -888
rect 1113 -936 1115 -932
rect 131 -950 213 -948
rect 247 -949 249 -946
rect 1129 -949 1131 -872
rect 1493 -871 1495 -865
rect 1493 -873 1513 -871
rect 1493 -885 1495 -882
rect 1156 -888 1158 -885
rect 1156 -946 1158 -928
rect 211 -972 213 -950
rect 105 -980 108 -978
rect 128 -980 146 -978
rect 186 -980 189 -978
rect 1113 -951 1131 -949
rect 1113 -957 1115 -951
rect 211 -995 213 -992
rect 131 -1002 213 -1000
rect 211 -1005 213 -1002
rect 247 -1007 249 -989
rect 1156 -969 1158 -966
rect 1493 -971 1495 -965
rect 1478 -973 1495 -971
rect 1478 -990 1480 -973
rect 1511 -990 1513 -873
rect 1744 -873 1746 -867
rect 1744 -875 1764 -873
rect 1744 -887 1746 -884
rect 1542 -922 1544 -919
rect 1542 -980 1544 -962
rect 1744 -973 1746 -967
rect 1729 -975 1746 -973
rect 1113 -1000 1115 -997
rect 211 -1028 213 -1025
rect 1729 -992 1731 -975
rect 1762 -992 1764 -875
rect 1793 -924 1795 -921
rect 1793 -982 1795 -964
rect 1542 -1003 1544 -1000
rect 1478 -1013 1480 -1010
rect 1511 -1013 1513 -1010
rect 2031 -993 2113 -991
rect 2147 -992 2149 -989
rect 1793 -1005 1795 -1002
rect 1729 -1015 1731 -1012
rect 1762 -1015 1764 -1012
rect 2111 -1015 2113 -993
rect 2005 -1023 2008 -1021
rect 2028 -1023 2046 -1021
rect 2086 -1023 2089 -1021
rect 105 -1031 108 -1029
rect 128 -1031 146 -1029
rect 186 -1031 189 -1029
rect 247 -1030 249 -1027
rect 2111 -1038 2113 -1035
rect 2031 -1045 2113 -1043
rect 2111 -1048 2113 -1045
rect 1017 -1063 1019 -1060
rect 1044 -1063 1046 -1060
rect 1235 -1063 1237 -1060
rect 1262 -1063 1264 -1060
rect 164 -1093 166 -1090
rect 191 -1093 193 -1090
rect 2147 -1050 2149 -1032
rect 2111 -1071 2113 -1068
rect 2005 -1074 2008 -1072
rect 2028 -1074 2046 -1072
rect 2086 -1074 2089 -1072
rect 2147 -1073 2149 -1070
rect 1017 -1131 1019 -1103
rect 1044 -1115 1046 -1103
rect 1044 -1117 1054 -1115
rect 1017 -1133 1038 -1131
rect -3284 -1156 -3282 -1153
rect -3556 -1184 -3474 -1182
rect -3440 -1183 -3438 -1180
rect -3476 -1206 -3474 -1184
rect -3582 -1214 -3579 -1212
rect -3559 -1214 -3541 -1212
rect -3501 -1214 -3498 -1212
rect -3349 -1199 -3347 -1196
rect -3476 -1229 -3474 -1226
rect -3556 -1236 -3474 -1234
rect -3476 -1239 -3474 -1236
rect -3440 -1241 -3438 -1223
rect 164 -1161 166 -1133
rect 191 -1145 193 -1133
rect 1036 -1137 1038 -1133
rect 191 -1147 201 -1145
rect 164 -1163 185 -1161
rect -3175 -1168 -3173 -1165
rect -3148 -1168 -3146 -1165
rect 183 -1167 185 -1163
rect -3476 -1262 -3474 -1259
rect -3349 -1257 -3347 -1239
rect -3284 -1242 -3282 -1236
rect -3175 -1236 -3173 -1208
rect -3148 -1220 -3146 -1208
rect 183 -1211 185 -1207
rect -3148 -1222 -3138 -1220
rect -3175 -1238 -3154 -1236
rect -3156 -1242 -3154 -1238
rect -3284 -1244 -3264 -1242
rect -3284 -1256 -3282 -1253
rect -3582 -1265 -3579 -1263
rect -3559 -1265 -3541 -1263
rect -3501 -1265 -3498 -1263
rect -3440 -1264 -3438 -1261
rect -3349 -1280 -3347 -1277
rect -3284 -1342 -3282 -1336
rect -3299 -1344 -3282 -1342
rect -3299 -1361 -3297 -1344
rect -3266 -1361 -3264 -1244
rect -3156 -1286 -3154 -1282
rect -3235 -1293 -3233 -1290
rect -3140 -1299 -3138 -1222
rect 199 -1224 201 -1147
rect 226 -1163 228 -1160
rect 1036 -1181 1038 -1177
rect 1052 -1194 1054 -1117
rect 1079 -1133 1081 -1130
rect 1235 -1131 1237 -1103
rect 1262 -1115 1264 -1103
rect 1262 -1117 1272 -1115
rect 1235 -1133 1256 -1131
rect 1254 -1137 1256 -1133
rect 1079 -1191 1081 -1173
rect 1254 -1181 1256 -1177
rect 1036 -1196 1054 -1194
rect 1036 -1202 1038 -1196
rect 226 -1221 228 -1203
rect 183 -1226 201 -1224
rect 183 -1232 185 -1226
rect -3113 -1238 -3111 -1235
rect 226 -1244 228 -1241
rect 1270 -1194 1272 -1117
rect 1297 -1133 1299 -1130
rect 1297 -1191 1299 -1173
rect 1254 -1196 1272 -1194
rect 1254 -1202 1256 -1196
rect 1079 -1214 1081 -1211
rect 1297 -1214 1299 -1211
rect 1036 -1245 1038 -1242
rect 1254 -1245 1256 -1242
rect 183 -1275 185 -1272
rect -3113 -1296 -3111 -1278
rect -3156 -1301 -3138 -1299
rect -3156 -1307 -3154 -1301
rect -3235 -1351 -3233 -1333
rect -3113 -1319 -3111 -1316
rect -3156 -1350 -3154 -1347
rect 779 -1355 781 -1352
rect 806 -1355 808 -1352
rect -3235 -1374 -3233 -1371
rect -3299 -1384 -3297 -1381
rect -3266 -1384 -3264 -1381
rect 779 -1423 781 -1395
rect 806 -1407 808 -1395
rect 806 -1409 816 -1407
rect 779 -1425 800 -1423
rect 798 -1429 800 -1425
rect 798 -1473 800 -1469
rect 814 -1486 816 -1409
rect 841 -1425 843 -1422
rect 841 -1483 843 -1465
rect 1430 -1482 1432 -1479
rect 798 -1488 816 -1486
rect 798 -1494 800 -1488
rect 841 -1506 843 -1503
rect 798 -1537 800 -1534
rect 1430 -1568 1432 -1562
rect 1430 -1570 1450 -1568
rect 1430 -1582 1432 -1579
rect 1016 -1585 1018 -1582
rect 1043 -1585 1045 -1582
rect 140 -1610 222 -1608
rect 256 -1609 258 -1606
rect 220 -1632 222 -1610
rect 114 -1640 117 -1638
rect 137 -1640 155 -1638
rect 195 -1640 198 -1638
rect 780 -1638 782 -1635
rect 807 -1638 809 -1635
rect 220 -1655 222 -1652
rect 140 -1662 222 -1660
rect 220 -1665 222 -1662
rect 256 -1667 258 -1649
rect 220 -1688 222 -1685
rect 1016 -1653 1018 -1625
rect 1043 -1637 1045 -1625
rect 1043 -1639 1053 -1637
rect 1016 -1655 1037 -1653
rect 1035 -1659 1037 -1655
rect 114 -1691 117 -1689
rect 137 -1691 155 -1689
rect 195 -1691 198 -1689
rect 256 -1690 258 -1687
rect 780 -1706 782 -1678
rect 807 -1690 809 -1678
rect 807 -1692 817 -1690
rect 780 -1708 801 -1706
rect 799 -1712 801 -1708
rect 173 -1753 175 -1750
rect 200 -1753 202 -1750
rect 799 -1756 801 -1752
rect 815 -1769 817 -1692
rect 1035 -1703 1037 -1699
rect 842 -1708 844 -1705
rect 1051 -1716 1053 -1639
rect 1078 -1655 1080 -1652
rect 1430 -1668 1432 -1662
rect 1415 -1670 1432 -1668
rect 1415 -1687 1417 -1670
rect 1448 -1687 1450 -1570
rect 1479 -1619 1481 -1616
rect 1727 -1635 1729 -1632
rect 1479 -1677 1481 -1659
rect 1078 -1713 1080 -1695
rect 1479 -1700 1481 -1697
rect 1415 -1710 1417 -1707
rect 1448 -1710 1450 -1707
rect 1035 -1718 1053 -1716
rect 1035 -1724 1037 -1718
rect 842 -1766 844 -1748
rect 2029 -1701 2111 -1699
rect 2145 -1700 2147 -1697
rect 1727 -1721 1729 -1715
rect 1727 -1723 1747 -1721
rect 2109 -1723 2111 -1701
rect 1078 -1736 1080 -1733
rect 1727 -1735 1729 -1732
rect 799 -1771 817 -1769
rect 799 -1777 801 -1771
rect 173 -1821 175 -1793
rect 200 -1805 202 -1793
rect 200 -1807 210 -1805
rect 173 -1823 194 -1821
rect 192 -1827 194 -1823
rect 192 -1871 194 -1867
rect 208 -1884 210 -1807
rect 1035 -1767 1037 -1764
rect 1441 -1782 1443 -1779
rect 842 -1789 844 -1786
rect 1025 -1796 1027 -1793
rect 1052 -1796 1054 -1793
rect 799 -1820 801 -1817
rect 235 -1823 237 -1820
rect 235 -1881 237 -1863
rect 1025 -1864 1027 -1836
rect 1052 -1848 1054 -1836
rect 1052 -1850 1062 -1848
rect 1025 -1866 1046 -1864
rect 1044 -1870 1046 -1866
rect 192 -1886 210 -1884
rect 192 -1892 194 -1886
rect 235 -1904 237 -1901
rect 776 -1909 778 -1906
rect 803 -1909 805 -1906
rect 192 -1935 194 -1932
rect 1044 -1914 1046 -1910
rect 1060 -1927 1062 -1850
rect 1727 -1821 1729 -1815
rect 1712 -1823 1729 -1821
rect 1712 -1840 1714 -1823
rect 1745 -1840 1747 -1723
rect 2003 -1731 2006 -1729
rect 2026 -1731 2044 -1729
rect 2084 -1731 2087 -1729
rect 2109 -1746 2111 -1743
rect 2029 -1753 2111 -1751
rect 2109 -1756 2111 -1753
rect 1776 -1772 1778 -1769
rect 2145 -1758 2147 -1740
rect 2109 -1779 2111 -1776
rect 2003 -1782 2006 -1780
rect 2026 -1782 2044 -1780
rect 2084 -1782 2087 -1780
rect 2145 -1781 2147 -1778
rect 1776 -1830 1778 -1812
rect 1776 -1853 1778 -1850
rect 1087 -1866 1089 -1863
rect 1441 -1868 1443 -1862
rect 1712 -1863 1714 -1860
rect 1745 -1863 1747 -1860
rect 1441 -1870 1461 -1868
rect 1441 -1882 1443 -1879
rect 1087 -1924 1089 -1906
rect 1044 -1929 1062 -1927
rect 1044 -1935 1046 -1929
rect 776 -1977 778 -1949
rect 803 -1961 805 -1949
rect 803 -1963 813 -1961
rect 776 -1979 797 -1977
rect 795 -1983 797 -1979
rect 795 -2027 797 -2023
rect 811 -2040 813 -1963
rect 1087 -1947 1089 -1944
rect 1441 -1968 1443 -1962
rect 1426 -1970 1443 -1968
rect 838 -1979 840 -1976
rect 1044 -1978 1046 -1975
rect 1426 -1987 1428 -1970
rect 1459 -1987 1461 -1870
rect 1490 -1919 1492 -1916
rect 1490 -1977 1492 -1959
rect 1490 -2000 1492 -1997
rect 1426 -2010 1428 -2007
rect 1459 -2010 1461 -2007
rect 838 -2037 840 -2019
rect 795 -2042 813 -2040
rect 795 -2048 797 -2042
rect 838 -2060 840 -2057
rect 795 -2091 797 -2088
rect 764 -2158 766 -2155
rect 791 -2158 793 -2155
rect 764 -2226 766 -2198
rect 791 -2210 793 -2198
rect 791 -2212 801 -2210
rect 764 -2228 785 -2226
rect 783 -2232 785 -2228
rect 783 -2276 785 -2272
rect 799 -2289 801 -2212
rect 826 -2228 828 -2225
rect 826 -2286 828 -2268
rect 783 -2291 801 -2289
rect 783 -2297 785 -2291
rect 826 -2309 828 -2306
rect 783 -2340 785 -2337
rect 137 -2485 219 -2483
rect 253 -2484 255 -2481
rect 217 -2507 219 -2485
rect 111 -2515 114 -2513
rect 134 -2515 152 -2513
rect 192 -2515 195 -2513
rect 1470 -2500 1472 -2497
rect 805 -2507 807 -2504
rect 832 -2507 834 -2504
rect 217 -2530 219 -2527
rect 137 -2537 219 -2535
rect 217 -2540 219 -2537
rect 253 -2542 255 -2524
rect 217 -2563 219 -2560
rect 111 -2566 114 -2564
rect 134 -2566 152 -2564
rect 192 -2566 195 -2564
rect 253 -2565 255 -2562
rect 805 -2575 807 -2547
rect 832 -2559 834 -2547
rect 1140 -2559 1142 -2556
rect 1167 -2559 1169 -2556
rect 832 -2561 842 -2559
rect 805 -2577 826 -2575
rect 824 -2581 826 -2577
rect 824 -2625 826 -2621
rect 170 -2628 172 -2625
rect 197 -2628 199 -2625
rect 840 -2638 842 -2561
rect 867 -2577 869 -2574
rect 2205 -2524 2207 -2521
rect 1470 -2586 1472 -2580
rect 1470 -2588 1490 -2586
rect 867 -2635 869 -2617
rect 1140 -2627 1142 -2599
rect 1167 -2611 1169 -2599
rect 1470 -2600 1472 -2597
rect 1167 -2613 1177 -2611
rect 1140 -2629 1161 -2627
rect 1159 -2633 1161 -2629
rect 824 -2640 842 -2638
rect 824 -2646 826 -2640
rect 170 -2696 172 -2668
rect 197 -2680 199 -2668
rect 197 -2682 207 -2680
rect 170 -2698 191 -2696
rect 189 -2702 191 -2698
rect 189 -2746 191 -2742
rect 205 -2759 207 -2682
rect 867 -2658 869 -2655
rect 1159 -2677 1161 -2673
rect 824 -2689 826 -2686
rect 1175 -2690 1177 -2613
rect 1202 -2629 1204 -2626
rect 1202 -2687 1204 -2669
rect 1470 -2686 1472 -2680
rect 232 -2698 234 -2695
rect 1159 -2692 1177 -2690
rect 1159 -2698 1161 -2692
rect 1455 -2688 1472 -2686
rect 1455 -2705 1457 -2688
rect 1488 -2705 1490 -2588
rect 2205 -2610 2207 -2604
rect 2205 -2612 2225 -2610
rect 2205 -2624 2207 -2621
rect 1519 -2637 1521 -2634
rect 1519 -2695 1521 -2677
rect 1202 -2710 1204 -2707
rect 2205 -2710 2207 -2704
rect 2190 -2712 2207 -2710
rect 1519 -2718 1521 -2715
rect 1455 -2728 1457 -2725
rect 1488 -2728 1490 -2725
rect 2190 -2729 2192 -2712
rect 2223 -2729 2225 -2612
rect 2254 -2661 2256 -2658
rect 2254 -2719 2256 -2701
rect 232 -2756 234 -2738
rect 1159 -2741 1161 -2738
rect 2254 -2742 2256 -2739
rect 2190 -2752 2192 -2749
rect 2223 -2752 2225 -2749
rect 189 -2761 207 -2759
rect 189 -2767 191 -2761
rect 232 -2779 234 -2776
rect 806 -2790 808 -2787
rect 833 -2790 835 -2787
rect 189 -2810 191 -2807
rect 806 -2858 808 -2830
rect 833 -2842 835 -2830
rect 1141 -2842 1143 -2839
rect 1168 -2842 1170 -2839
rect 833 -2844 843 -2842
rect 806 -2860 827 -2858
rect 825 -2864 827 -2860
rect 825 -2908 827 -2904
rect 841 -2921 843 -2844
rect 868 -2860 870 -2857
rect 868 -2918 870 -2900
rect 1141 -2910 1143 -2882
rect 1168 -2894 1170 -2882
rect 1477 -2889 1479 -2886
rect 1168 -2896 1178 -2894
rect 1141 -2912 1162 -2910
rect 1160 -2916 1162 -2912
rect 825 -2923 843 -2921
rect 825 -2929 827 -2923
rect 868 -2941 870 -2938
rect 1160 -2960 1162 -2956
rect 825 -2972 827 -2969
rect 1176 -2973 1178 -2896
rect 1203 -2912 1205 -2909
rect 1203 -2970 1205 -2952
rect 1160 -2975 1178 -2973
rect 1160 -2981 1162 -2975
rect 1477 -2975 1479 -2969
rect 1477 -2977 1497 -2975
rect 1477 -2989 1479 -2986
rect 1203 -2993 1205 -2990
rect 1160 -3024 1162 -3021
rect 802 -3061 804 -3058
rect 829 -3061 831 -3058
rect 1477 -3075 1479 -3069
rect 1462 -3077 1479 -3075
rect 1462 -3094 1464 -3077
rect 1495 -3094 1497 -2977
rect 1526 -3026 1528 -3023
rect 1769 -3045 1771 -3042
rect 1526 -3084 1528 -3066
rect 802 -3129 804 -3101
rect 829 -3113 831 -3101
rect 829 -3115 839 -3113
rect 1526 -3107 1528 -3104
rect 802 -3131 823 -3129
rect 821 -3135 823 -3131
rect 821 -3179 823 -3175
rect 837 -3192 839 -3115
rect 1462 -3117 1464 -3114
rect 1495 -3117 1497 -3114
rect 864 -3131 866 -3128
rect 1769 -3131 1771 -3125
rect 1769 -3133 1789 -3131
rect 1769 -3145 1771 -3142
rect 864 -3189 866 -3171
rect 821 -3194 839 -3192
rect 821 -3200 823 -3194
rect 864 -3212 866 -3209
rect 1769 -3231 1771 -3225
rect 1754 -3233 1771 -3231
rect 821 -3243 823 -3240
rect 1471 -3244 1473 -3241
rect 1498 -3244 1500 -3241
rect 1754 -3250 1756 -3233
rect 1787 -3250 1789 -3133
rect 1818 -3182 1820 -3179
rect 1818 -3240 1820 -3222
rect 1818 -3263 1820 -3260
rect 1754 -3273 1756 -3270
rect 1787 -3273 1789 -3270
rect 790 -3310 792 -3307
rect 817 -3310 819 -3307
rect 1471 -3312 1473 -3284
rect 1498 -3296 1500 -3284
rect 1498 -3298 1508 -3296
rect 1471 -3314 1492 -3312
rect 1490 -3318 1492 -3314
rect 790 -3378 792 -3350
rect 817 -3362 819 -3350
rect 1490 -3362 1492 -3358
rect 817 -3364 827 -3362
rect 790 -3380 811 -3378
rect 809 -3384 811 -3380
rect 809 -3428 811 -3424
rect 825 -3441 827 -3364
rect 1131 -3376 1133 -3373
rect 1158 -3376 1160 -3373
rect 1506 -3375 1508 -3298
rect 1533 -3314 1535 -3311
rect 1533 -3372 1535 -3354
rect 852 -3380 854 -3377
rect 1490 -3377 1508 -3375
rect 1490 -3383 1492 -3377
rect 852 -3438 854 -3420
rect 809 -3443 827 -3441
rect 809 -3449 811 -3443
rect 1131 -3444 1133 -3416
rect 1158 -3428 1160 -3416
rect 1533 -3395 1535 -3392
rect 1490 -3426 1492 -3423
rect 1158 -3430 1168 -3428
rect 1131 -3446 1152 -3444
rect 1150 -3450 1152 -3446
rect 852 -3461 854 -3458
rect 809 -3492 811 -3489
rect 1150 -3494 1152 -3490
rect 1166 -3507 1168 -3430
rect 1193 -3446 1195 -3443
rect 1193 -3504 1195 -3486
rect 1150 -3509 1168 -3507
rect 1150 -3515 1152 -3509
rect 1193 -3527 1195 -3524
rect 1150 -3558 1152 -3555
rect 807 -3577 809 -3574
rect 834 -3577 836 -3574
rect 807 -3645 809 -3617
rect 834 -3629 836 -3617
rect 834 -3631 844 -3629
rect 807 -3647 828 -3645
rect 826 -3651 828 -3647
rect 826 -3695 828 -3691
rect 842 -3708 844 -3631
rect 869 -3647 871 -3644
rect 869 -3705 871 -3687
rect 826 -3710 844 -3708
rect 826 -3716 828 -3710
rect 869 -3728 871 -3725
rect 826 -3759 828 -3756
rect 795 -3826 797 -3823
rect 822 -3826 824 -3823
rect 795 -3894 797 -3866
rect 822 -3878 824 -3866
rect 822 -3880 832 -3878
rect 795 -3896 816 -3894
rect 814 -3900 816 -3896
rect 814 -3944 816 -3940
rect 830 -3957 832 -3880
rect 857 -3896 859 -3893
rect 857 -3954 859 -3936
rect 814 -3959 832 -3957
rect 814 -3965 816 -3959
rect 857 -3977 859 -3974
rect 814 -4008 816 -4005
<< polycontact >>
rect 1619 32 1624 37
rect 1619 9 1624 14
rect 1619 -13 1624 -8
rect 1730 -17 1735 -12
rect 1619 -42 1624 -37
rect 143 -169 148 -164
rect 143 -192 148 -187
rect 1099 -151 1104 -146
rect 143 -214 148 -209
rect 254 -218 259 -213
rect 143 -243 148 -238
rect 729 -218 734 -213
rect 1084 -254 1089 -249
rect 791 -273 796 -268
rect 1614 -188 1619 -183
rect 1614 -211 1619 -206
rect 1614 -233 1619 -228
rect 1725 -237 1730 -232
rect 1148 -255 1153 -250
rect 748 -284 753 -279
rect 1614 -262 1619 -257
rect 171 -377 176 -372
rect 233 -432 238 -427
rect 190 -443 195 -438
rect 1089 -888 1094 -883
rect 1488 -873 1493 -868
rect 1151 -943 1156 -938
rect 131 -955 136 -950
rect 131 -978 136 -973
rect 1108 -954 1113 -949
rect 131 -1000 136 -995
rect 242 -1004 247 -999
rect 131 -1029 136 -1024
rect 1473 -976 1478 -971
rect 1739 -875 1744 -870
rect 1537 -977 1542 -972
rect 1724 -978 1729 -973
rect 1788 -979 1793 -974
rect 2031 -998 2036 -993
rect 2031 -1021 2036 -1016
rect 2031 -1043 2036 -1038
rect 2142 -1047 2147 -1042
rect 2031 -1072 2036 -1067
rect 1012 -1133 1017 -1128
rect -3556 -1189 -3551 -1184
rect -3556 -1212 -3551 -1207
rect -3556 -1234 -3551 -1229
rect -3445 -1238 -3440 -1233
rect -3556 -1263 -3551 -1258
rect 159 -1163 164 -1158
rect -3354 -1254 -3349 -1249
rect -3289 -1244 -3284 -1239
rect -3180 -1238 -3175 -1233
rect -3304 -1347 -3299 -1342
rect 1230 -1133 1235 -1128
rect 1074 -1188 1079 -1183
rect 1031 -1199 1036 -1194
rect 221 -1218 226 -1213
rect 178 -1229 183 -1224
rect 1292 -1188 1297 -1183
rect 1249 -1199 1254 -1194
rect -3118 -1293 -3113 -1288
rect -3161 -1304 -3156 -1299
rect -3240 -1348 -3235 -1343
rect 774 -1425 779 -1420
rect 836 -1480 841 -1475
rect 793 -1491 798 -1486
rect 1425 -1570 1430 -1565
rect 140 -1615 145 -1610
rect 140 -1638 145 -1633
rect 140 -1660 145 -1655
rect 251 -1664 256 -1659
rect 140 -1689 145 -1684
rect 1011 -1655 1016 -1650
rect 775 -1708 780 -1703
rect 1410 -1673 1415 -1668
rect 1474 -1674 1479 -1669
rect 1073 -1710 1078 -1705
rect 1030 -1721 1035 -1716
rect 837 -1763 842 -1758
rect 2029 -1706 2034 -1701
rect 1722 -1723 1727 -1718
rect 794 -1774 799 -1769
rect 168 -1823 173 -1818
rect 230 -1878 235 -1873
rect 1020 -1866 1025 -1861
rect 187 -1889 192 -1884
rect 1707 -1826 1712 -1821
rect 2029 -1729 2034 -1724
rect 2029 -1751 2034 -1746
rect 2140 -1755 2145 -1750
rect 2029 -1780 2034 -1775
rect 1771 -1827 1776 -1822
rect 1436 -1870 1441 -1865
rect 1082 -1921 1087 -1916
rect 1039 -1932 1044 -1927
rect 771 -1979 776 -1974
rect 1421 -1973 1426 -1968
rect 1485 -1974 1490 -1969
rect 833 -2034 838 -2029
rect 790 -2045 795 -2040
rect 759 -2228 764 -2223
rect 821 -2283 826 -2278
rect 778 -2294 783 -2289
rect 137 -2490 142 -2485
rect 137 -2513 142 -2508
rect 137 -2535 142 -2530
rect 248 -2539 253 -2534
rect 137 -2564 142 -2559
rect 800 -2577 805 -2572
rect 1465 -2588 1470 -2583
rect 862 -2632 867 -2627
rect 1135 -2629 1140 -2624
rect 819 -2643 824 -2638
rect 165 -2698 170 -2693
rect 1197 -2684 1202 -2679
rect 1154 -2695 1159 -2690
rect 1450 -2691 1455 -2686
rect 2200 -2612 2205 -2607
rect 1514 -2692 1519 -2687
rect 2185 -2715 2190 -2710
rect 2249 -2716 2254 -2711
rect 227 -2753 232 -2748
rect 184 -2764 189 -2759
rect 801 -2860 806 -2855
rect 863 -2915 868 -2910
rect 1136 -2912 1141 -2907
rect 820 -2926 825 -2921
rect 1198 -2967 1203 -2962
rect 1155 -2978 1160 -2973
rect 1472 -2977 1477 -2972
rect 1457 -3080 1462 -3075
rect 1521 -3081 1526 -3076
rect 797 -3131 802 -3126
rect 1764 -3133 1769 -3128
rect 859 -3186 864 -3181
rect 816 -3197 821 -3192
rect 1749 -3236 1754 -3231
rect 1813 -3237 1818 -3232
rect 1466 -3314 1471 -3309
rect 785 -3380 790 -3375
rect 1528 -3369 1533 -3364
rect 1485 -3380 1490 -3375
rect 847 -3435 852 -3430
rect 804 -3446 809 -3441
rect 1126 -3446 1131 -3441
rect 1188 -3501 1193 -3496
rect 1145 -3512 1150 -3507
rect 802 -3647 807 -3642
rect 864 -3702 869 -3697
rect 821 -3713 826 -3708
rect 790 -3896 795 -3891
rect 852 -3951 857 -3946
rect 809 -3962 814 -3957
<< metal1 >>
rect 1722 49 1749 52
rect 1722 45 1725 49
rect 1729 45 1742 49
rect 1746 45 1749 49
rect 1722 43 1749 45
rect 1730 38 1734 43
rect -31 26 299 30
rect 1619 30 1624 32
rect 304 26 1624 30
rect 741 25 1624 26
rect 1584 21 1590 22
rect 1584 17 1585 21
rect 1589 17 1590 21
rect 1584 14 1590 17
rect 1619 14 1624 25
rect 1679 19 1688 22
rect 1679 15 1681 19
rect 1685 15 1688 19
rect 1702 15 1715 18
rect 1679 14 1688 15
rect 1584 10 1596 14
rect 1584 0 1590 10
rect 1674 10 1688 14
rect 1616 2 1634 6
rect 1679 2 1688 10
rect 1584 -4 1585 0
rect 1589 -4 1590 0
rect 1584 -5 1590 -4
rect 1619 -8 1624 2
rect 1679 -2 1681 2
rect 1685 -2 1688 2
rect 1679 -5 1688 -2
rect 1694 -8 1698 -5
rect 1648 -12 1698 -8
rect 1648 -17 1652 -12
rect 313 -22 1652 -17
rect 1702 -18 1706 -5
rect 1709 -12 1715 15
rect 1738 -12 1742 -2
rect 1709 -17 1730 -12
rect 1738 -17 1787 -12
rect 1584 -30 1590 -29
rect 1584 -34 1585 -30
rect 1589 -34 1590 -30
rect 1584 -37 1590 -34
rect 1619 -37 1624 -22
rect 1679 -32 1688 -29
rect 1679 -36 1681 -32
rect 1685 -36 1688 -32
rect 1679 -37 1688 -36
rect 1584 -41 1596 -37
rect 1091 -52 1118 -49
rect 1091 -56 1094 -52
rect 1098 -56 1111 -52
rect 1115 -56 1118 -52
rect 1584 -51 1590 -41
rect 1674 -41 1688 -37
rect 1616 -49 1634 -45
rect 1679 -49 1688 -41
rect 1584 -55 1585 -51
rect 1589 -55 1590 -51
rect 1584 -56 1590 -55
rect 1091 -58 1118 -56
rect 1099 -63 1103 -58
rect 721 -137 775 -134
rect 721 -141 724 -137
rect 728 -141 741 -137
rect 745 -141 751 -137
rect 755 -141 768 -137
rect 772 -141 775 -137
rect 721 -143 775 -141
rect 1619 -69 1624 -49
rect 1679 -53 1681 -49
rect 1685 -53 1688 -49
rect 1679 -56 1688 -53
rect 1738 -20 1742 -17
rect 1694 -69 1698 -38
rect 1730 -46 1734 -40
rect 1722 -47 1749 -46
rect 1722 -51 1723 -47
rect 1727 -51 1744 -47
rect 1748 -51 1749 -47
rect 1722 -52 1749 -51
rect 1619 -72 1698 -69
rect 729 -148 733 -143
rect 756 -148 760 -143
rect 246 -152 273 -149
rect 246 -156 249 -152
rect 253 -156 266 -152
rect 270 -156 273 -152
rect 246 -158 273 -156
rect 254 -163 258 -158
rect 143 -171 148 -169
rect -19 -176 14 -171
rect 19 -176 148 -171
rect 108 -180 114 -179
rect 108 -184 109 -180
rect 113 -184 114 -180
rect 108 -187 114 -184
rect 143 -187 148 -176
rect 203 -182 212 -179
rect 203 -186 205 -182
rect 209 -186 212 -182
rect 226 -186 239 -183
rect 203 -187 212 -186
rect 108 -191 120 -187
rect 108 -201 114 -191
rect 198 -191 212 -187
rect 140 -199 158 -195
rect 203 -199 212 -191
rect 108 -205 109 -201
rect 113 -205 114 -201
rect 108 -206 114 -205
rect 143 -209 148 -199
rect 203 -203 205 -199
rect 209 -203 212 -199
rect 203 -206 212 -203
rect 218 -209 222 -206
rect 172 -213 222 -209
rect 172 -218 176 -213
rect -16 -223 176 -218
rect 226 -219 230 -206
rect 233 -213 239 -186
rect 262 -213 266 -203
rect 737 -208 741 -188
rect 764 -208 768 -188
rect 1011 -151 1099 -146
rect 783 -207 810 -204
rect 737 -212 778 -208
rect 233 -218 254 -213
rect 262 -218 308 -213
rect 313 -218 729 -213
rect 69 -438 74 -223
rect 108 -231 114 -230
rect 108 -235 109 -231
rect 113 -235 114 -231
rect 108 -238 114 -235
rect 143 -238 148 -223
rect 203 -233 212 -230
rect 203 -237 205 -233
rect 209 -237 212 -233
rect 203 -238 212 -237
rect 108 -242 120 -238
rect 108 -252 114 -242
rect 198 -242 212 -238
rect 140 -250 158 -246
rect 203 -250 212 -242
rect 108 -256 109 -252
rect 113 -256 114 -252
rect 108 -257 114 -256
rect 143 -270 148 -250
rect 203 -254 205 -250
rect 209 -254 212 -250
rect 203 -257 212 -254
rect 262 -221 266 -218
rect 218 -270 222 -239
rect 756 -222 760 -212
rect 254 -247 258 -241
rect 246 -248 273 -247
rect 246 -252 247 -248
rect 251 -252 268 -248
rect 272 -252 273 -248
rect 246 -253 273 -252
rect 143 -273 222 -270
rect 748 -268 752 -262
rect 773 -268 778 -212
rect 783 -211 786 -207
rect 790 -211 803 -207
rect 807 -211 810 -207
rect 783 -213 810 -211
rect 791 -218 795 -213
rect 799 -268 803 -258
rect 1011 -268 1016 -151
rect 1107 -155 1111 -143
rect 1099 -159 1111 -155
rect 1099 -163 1103 -159
rect 1717 -171 1744 -168
rect 1717 -175 1720 -171
rect 1724 -175 1737 -171
rect 1741 -175 1744 -171
rect 1717 -177 1744 -175
rect 1725 -182 1729 -177
rect 1140 -189 1167 -186
rect 1140 -193 1143 -189
rect 1147 -193 1160 -189
rect 1164 -193 1167 -189
rect 1614 -190 1619 -188
rect 1140 -195 1167 -193
rect 1542 -195 1619 -190
rect 1148 -200 1152 -195
rect 748 -272 762 -268
rect 756 -273 762 -272
rect 773 -273 791 -268
rect 799 -273 1016 -268
rect 1040 -254 1084 -249
rect 1107 -250 1111 -243
rect 1156 -250 1160 -240
rect 1542 -250 1547 -195
rect 1579 -199 1585 -198
rect 1579 -203 1580 -199
rect 1584 -203 1585 -199
rect 1579 -206 1585 -203
rect 1614 -206 1619 -195
rect 1674 -201 1683 -198
rect 1674 -205 1676 -201
rect 1680 -205 1683 -201
rect 1697 -205 1710 -202
rect 1674 -206 1683 -205
rect 1579 -210 1591 -206
rect 1579 -220 1585 -210
rect 1669 -210 1683 -206
rect 1611 -218 1629 -214
rect 1674 -218 1683 -210
rect 1579 -224 1580 -220
rect 1584 -224 1585 -220
rect 1579 -225 1585 -224
rect 1614 -228 1619 -218
rect 1674 -222 1676 -218
rect 1680 -222 1683 -218
rect 1674 -225 1683 -222
rect 1689 -228 1693 -225
rect 1643 -232 1693 -228
rect 1643 -237 1647 -232
rect 304 -284 748 -279
rect 756 -287 760 -273
rect 799 -276 803 -273
rect 163 -296 217 -293
rect 163 -300 166 -296
rect 170 -300 183 -296
rect 187 -300 193 -296
rect 197 -300 210 -296
rect 214 -300 217 -296
rect 163 -302 217 -300
rect 171 -307 175 -302
rect 198 -307 202 -302
rect 791 -302 795 -296
rect 783 -303 810 -302
rect 783 -307 784 -303
rect 788 -307 805 -303
rect 809 -307 810 -303
rect 783 -308 810 -307
rect 748 -333 752 -327
rect 740 -334 767 -333
rect 740 -338 741 -334
rect 745 -338 762 -334
rect 766 -338 767 -334
rect 740 -339 767 -338
rect 179 -367 183 -347
rect 206 -367 210 -347
rect 225 -366 252 -363
rect 179 -371 220 -367
rect 107 -377 171 -372
rect 198 -381 202 -371
rect 190 -427 194 -421
rect 215 -427 220 -371
rect 225 -370 228 -366
rect 232 -370 245 -366
rect 249 -370 252 -366
rect 225 -372 252 -370
rect 233 -377 237 -372
rect 241 -427 245 -417
rect 1040 -427 1045 -254
rect 1107 -255 1148 -250
rect 1156 -255 1547 -250
rect 1556 -242 1647 -237
rect 1697 -238 1701 -225
rect 1704 -232 1710 -205
rect 1733 -232 1737 -222
rect 1704 -237 1725 -232
rect 1733 -237 1789 -232
rect 1107 -258 1111 -255
rect 1156 -258 1160 -255
rect 1092 -262 1129 -258
rect 1092 -268 1096 -262
rect 1125 -268 1129 -262
rect 1148 -284 1152 -278
rect 1140 -285 1167 -284
rect 1084 -294 1088 -288
rect 1117 -294 1121 -288
rect 1140 -289 1141 -285
rect 1145 -289 1162 -285
rect 1166 -289 1167 -285
rect 1140 -290 1167 -289
rect 1076 -295 1103 -294
rect 1076 -299 1077 -295
rect 1081 -299 1098 -295
rect 1102 -299 1103 -295
rect 1076 -300 1103 -299
rect 1109 -295 1136 -294
rect 1109 -299 1110 -295
rect 1114 -299 1131 -295
rect 1135 -299 1136 -295
rect 1109 -300 1136 -299
rect 190 -431 204 -427
rect 198 -432 204 -431
rect 215 -432 233 -427
rect 241 -432 317 -427
rect 322 -432 1045 -427
rect 69 -443 190 -438
rect 198 -446 202 -432
rect 241 -435 245 -432
rect 233 -461 237 -455
rect 1556 -456 1561 -242
rect 1579 -250 1585 -249
rect 1579 -254 1580 -250
rect 1584 -254 1585 -250
rect 1579 -257 1585 -254
rect 1614 -257 1619 -242
rect 1674 -252 1683 -249
rect 1674 -256 1676 -252
rect 1680 -256 1683 -252
rect 1674 -257 1683 -256
rect 1579 -261 1591 -257
rect 1579 -271 1585 -261
rect 1669 -261 1683 -257
rect 1611 -269 1629 -265
rect 1674 -269 1683 -261
rect 1579 -275 1580 -271
rect 1584 -275 1585 -271
rect 1579 -276 1585 -275
rect 1614 -289 1619 -269
rect 1674 -273 1676 -269
rect 1680 -273 1683 -269
rect 1674 -276 1683 -273
rect 1733 -240 1737 -237
rect 1689 -289 1693 -258
rect 1725 -266 1729 -260
rect 1717 -267 1744 -266
rect 1717 -271 1718 -267
rect 1722 -271 1739 -267
rect 1743 -271 1744 -267
rect 1717 -272 1744 -271
rect 1614 -292 1693 -289
rect 331 -461 1561 -456
rect 225 -462 252 -461
rect 225 -466 226 -462
rect 230 -466 247 -462
rect 251 -466 252 -462
rect 225 -467 252 -466
rect 190 -492 194 -486
rect 182 -493 209 -492
rect 182 -497 183 -493
rect 187 -497 204 -493
rect 208 -497 209 -493
rect 182 -498 209 -497
rect 335 -757 1443 -752
rect 335 -859 340 -757
rect 1081 -807 1135 -804
rect 1081 -811 1084 -807
rect 1088 -811 1101 -807
rect 1105 -811 1111 -807
rect 1115 -811 1128 -807
rect 1132 -811 1135 -807
rect 1081 -813 1135 -811
rect 1089 -818 1093 -813
rect 1116 -818 1120 -813
rect 335 -867 340 -864
rect 1097 -878 1101 -858
rect 1124 -878 1128 -858
rect 1438 -868 1443 -757
rect 1480 -774 1507 -771
rect 1480 -778 1483 -774
rect 1487 -778 1500 -774
rect 1504 -778 1507 -774
rect 1480 -780 1507 -778
rect 1731 -776 1758 -773
rect 1731 -780 1734 -776
rect 1738 -780 1751 -776
rect 1755 -780 1758 -776
rect 1488 -785 1492 -780
rect 1731 -782 1758 -780
rect 1438 -873 1488 -868
rect 1143 -877 1170 -874
rect 1496 -877 1500 -865
rect 1739 -787 1743 -782
rect 1097 -882 1138 -878
rect 322 -888 1089 -883
rect 1116 -892 1120 -882
rect 234 -938 261 -935
rect 234 -942 237 -938
rect 241 -942 254 -938
rect 258 -942 261 -938
rect 1108 -938 1112 -932
rect 1133 -938 1138 -882
rect 1143 -881 1146 -877
rect 1150 -881 1163 -877
rect 1167 -881 1170 -877
rect 1143 -883 1170 -881
rect 1488 -881 1500 -877
rect 1660 -875 1739 -870
rect 1151 -888 1155 -883
rect 1488 -885 1492 -881
rect 1159 -938 1163 -928
rect 1108 -942 1122 -938
rect 234 -944 261 -942
rect 1116 -943 1122 -942
rect 1133 -943 1151 -938
rect 1159 -943 1466 -938
rect 242 -949 246 -944
rect 131 -957 136 -955
rect -31 -962 2 -957
rect 7 -962 136 -957
rect 96 -966 102 -965
rect 96 -970 97 -966
rect 101 -970 102 -966
rect 96 -973 102 -970
rect 131 -973 136 -962
rect 191 -968 200 -965
rect 191 -972 193 -968
rect 197 -972 200 -968
rect 214 -972 227 -969
rect 191 -973 200 -972
rect 96 -977 108 -973
rect 96 -987 102 -977
rect 186 -977 200 -973
rect 128 -985 146 -981
rect 191 -985 200 -977
rect 96 -991 97 -987
rect 101 -991 102 -987
rect 96 -992 102 -991
rect 131 -995 136 -985
rect 191 -989 193 -985
rect 197 -989 200 -985
rect 191 -992 200 -989
rect 206 -995 210 -992
rect 160 -999 210 -995
rect 160 -1004 164 -999
rect -28 -1009 164 -1004
rect 214 -1005 218 -992
rect 221 -999 227 -972
rect 250 -999 254 -989
rect 1043 -954 1108 -949
rect 1043 -999 1048 -954
rect 1116 -957 1120 -943
rect 1159 -946 1163 -943
rect 221 -1004 242 -999
rect 250 -1004 326 -999
rect 331 -1004 1048 -999
rect 1151 -972 1155 -966
rect 1461 -971 1466 -943
rect 1529 -911 1556 -908
rect 1529 -915 1532 -911
rect 1536 -915 1549 -911
rect 1553 -915 1556 -911
rect 1529 -917 1556 -915
rect 1537 -922 1541 -917
rect 1143 -973 1170 -972
rect 1143 -977 1144 -973
rect 1148 -977 1165 -973
rect 1169 -977 1170 -973
rect 1461 -976 1473 -971
rect 1496 -972 1500 -965
rect 1545 -972 1549 -962
rect 1660 -972 1665 -875
rect 1747 -879 1751 -867
rect 1739 -883 1751 -879
rect 1739 -887 1743 -883
rect 1780 -913 1807 -910
rect 1780 -917 1783 -913
rect 1787 -917 1800 -913
rect 1804 -917 1807 -913
rect 1780 -919 1807 -917
rect 1788 -924 1792 -919
rect 1143 -978 1170 -977
rect 1496 -977 1537 -972
rect 1545 -977 1665 -972
rect 1496 -980 1500 -977
rect 1545 -980 1549 -977
rect 1481 -984 1518 -980
rect 1481 -990 1485 -984
rect 1514 -990 1518 -984
rect 1108 -1003 1112 -997
rect 1100 -1004 1127 -1003
rect -3297 -1145 -3270 -1142
rect -3297 -1149 -3294 -1145
rect -3290 -1149 -3277 -1145
rect -3273 -1149 -3270 -1145
rect -3297 -1151 -3270 -1149
rect -3289 -1156 -3285 -1151
rect -3453 -1172 -3426 -1169
rect -3453 -1176 -3450 -1172
rect -3446 -1176 -3433 -1172
rect -3429 -1176 -3426 -1172
rect -3453 -1178 -3426 -1176
rect -3445 -1183 -3441 -1178
rect -3556 -1191 -3551 -1189
rect -3591 -1196 -3551 -1191
rect -3591 -1200 -3585 -1199
rect -3591 -1204 -3590 -1200
rect -3586 -1204 -3585 -1200
rect -3591 -1207 -3585 -1204
rect -3556 -1207 -3551 -1196
rect -3496 -1202 -3487 -1199
rect -3496 -1206 -3494 -1202
rect -3490 -1206 -3487 -1202
rect -3473 -1206 -3460 -1203
rect -3496 -1207 -3487 -1206
rect -3591 -1211 -3579 -1207
rect -3591 -1221 -3585 -1211
rect -3501 -1211 -3487 -1207
rect -3559 -1219 -3541 -1215
rect -3496 -1219 -3487 -1211
rect -3591 -1225 -3590 -1221
rect -3586 -1225 -3585 -1221
rect -3591 -1226 -3585 -1225
rect -3556 -1229 -3551 -1219
rect -3496 -1223 -3494 -1219
rect -3490 -1223 -3487 -1219
rect -3496 -1226 -3487 -1223
rect -3481 -1229 -3477 -1226
rect -3527 -1233 -3477 -1229
rect -3527 -1238 -3523 -1233
rect -3591 -1243 -3523 -1238
rect -3473 -1239 -3469 -1226
rect -3466 -1233 -3460 -1206
rect -3362 -1188 -3335 -1185
rect -3362 -1192 -3359 -1188
rect -3355 -1192 -3342 -1188
rect -3338 -1192 -3335 -1188
rect -3362 -1194 -3335 -1192
rect -3437 -1233 -3433 -1223
rect -3354 -1199 -3350 -1194
rect -3466 -1238 -3445 -1233
rect -3437 -1238 -3426 -1233
rect -3591 -1251 -3585 -1250
rect -3591 -1255 -3590 -1251
rect -3586 -1255 -3585 -1251
rect -3591 -1258 -3585 -1255
rect -3556 -1258 -3551 -1243
rect -3496 -1253 -3487 -1250
rect -3496 -1257 -3494 -1253
rect -3490 -1257 -3487 -1253
rect -3496 -1258 -3487 -1257
rect -3591 -1262 -3579 -1258
rect -3591 -1272 -3585 -1262
rect -3501 -1262 -3487 -1258
rect -3559 -1270 -3541 -1266
rect -3496 -1270 -3487 -1262
rect -3591 -1276 -3590 -1272
rect -3586 -1276 -3585 -1272
rect -3591 -1277 -3585 -1276
rect -3556 -1290 -3551 -1270
rect -3496 -1274 -3494 -1270
rect -3490 -1274 -3487 -1270
rect -3496 -1277 -3487 -1274
rect -3437 -1241 -3433 -1238
rect -3188 -1157 -3134 -1154
rect -3188 -1161 -3185 -1157
rect -3181 -1161 -3168 -1157
rect -3164 -1161 -3158 -1157
rect -3154 -1161 -3141 -1157
rect -3137 -1161 -3134 -1157
rect -3188 -1163 -3134 -1161
rect -3180 -1168 -3176 -1163
rect -3153 -1168 -3149 -1163
rect -3172 -1228 -3168 -1208
rect -3145 -1228 -3141 -1208
rect 57 -1224 62 -1009
rect 96 -1017 102 -1016
rect 96 -1021 97 -1017
rect 101 -1021 102 -1017
rect 96 -1024 102 -1021
rect 131 -1024 136 -1009
rect 191 -1019 200 -1016
rect 191 -1023 193 -1019
rect 197 -1023 200 -1019
rect 191 -1024 200 -1023
rect 96 -1028 108 -1024
rect 96 -1038 102 -1028
rect 186 -1028 200 -1024
rect 128 -1036 146 -1032
rect 191 -1036 200 -1028
rect 96 -1042 97 -1038
rect 101 -1042 102 -1038
rect 96 -1043 102 -1042
rect 131 -1056 136 -1036
rect 191 -1040 193 -1036
rect 197 -1040 200 -1036
rect 191 -1043 200 -1040
rect 250 -1007 254 -1004
rect 206 -1056 210 -1025
rect 1100 -1008 1101 -1004
rect 1105 -1008 1122 -1004
rect 1126 -1008 1127 -1004
rect 1100 -1009 1127 -1008
rect 1691 -978 1724 -973
rect 1747 -974 1751 -967
rect 1796 -974 1800 -964
rect 1537 -1006 1541 -1000
rect 1529 -1007 1556 -1006
rect 1473 -1016 1477 -1010
rect 1506 -1016 1510 -1010
rect 1529 -1011 1530 -1007
rect 1534 -1011 1551 -1007
rect 1555 -1011 1556 -1007
rect 1529 -1012 1556 -1011
rect 1465 -1017 1492 -1016
rect 1465 -1021 1466 -1017
rect 1470 -1021 1487 -1017
rect 1491 -1021 1492 -1017
rect 1465 -1022 1492 -1021
rect 1498 -1017 1525 -1016
rect 1498 -1021 1499 -1017
rect 1503 -1021 1520 -1017
rect 1524 -1021 1525 -1017
rect 1498 -1022 1525 -1021
rect 242 -1033 246 -1027
rect 234 -1034 261 -1033
rect 234 -1038 235 -1034
rect 239 -1038 256 -1034
rect 260 -1038 261 -1034
rect 234 -1039 261 -1038
rect 131 -1059 210 -1056
rect 1004 -1052 1058 -1049
rect 1004 -1056 1007 -1052
rect 1011 -1056 1024 -1052
rect 1028 -1056 1034 -1052
rect 1038 -1056 1051 -1052
rect 1055 -1056 1058 -1052
rect 1004 -1058 1058 -1056
rect 1222 -1052 1276 -1049
rect 1222 -1056 1225 -1052
rect 1229 -1056 1242 -1052
rect 1246 -1056 1252 -1052
rect 1256 -1056 1269 -1052
rect 1273 -1056 1276 -1052
rect 1222 -1058 1276 -1056
rect 1012 -1063 1016 -1058
rect 1039 -1063 1043 -1058
rect 1230 -1063 1234 -1058
rect 1257 -1063 1261 -1058
rect 151 -1082 205 -1079
rect 151 -1086 154 -1082
rect 158 -1086 171 -1082
rect 175 -1086 181 -1082
rect 185 -1086 198 -1082
rect 202 -1086 205 -1082
rect 151 -1088 205 -1086
rect 159 -1093 163 -1088
rect 186 -1093 190 -1088
rect 1020 -1123 1024 -1103
rect 1047 -1123 1051 -1103
rect 1066 -1122 1093 -1119
rect 1020 -1127 1061 -1123
rect 304 -1133 1012 -1128
rect 167 -1153 171 -1133
rect 194 -1153 198 -1133
rect 1039 -1137 1043 -1127
rect 313 -1145 1000 -1140
rect 213 -1152 240 -1149
rect 167 -1157 208 -1153
rect 95 -1163 159 -1158
rect 186 -1167 190 -1157
rect 178 -1213 182 -1207
rect 203 -1213 208 -1157
rect 213 -1156 216 -1152
rect 220 -1156 233 -1152
rect 237 -1156 240 -1152
rect 213 -1158 240 -1156
rect 221 -1163 225 -1158
rect 995 -1194 1000 -1145
rect 1031 -1183 1035 -1177
rect 1056 -1183 1061 -1127
rect 1066 -1126 1069 -1122
rect 1073 -1126 1086 -1122
rect 1090 -1126 1093 -1122
rect 1066 -1128 1093 -1126
rect 1238 -1123 1242 -1103
rect 1265 -1123 1269 -1103
rect 1284 -1122 1311 -1119
rect 1238 -1127 1279 -1123
rect 1186 -1128 1218 -1127
rect 1074 -1133 1078 -1128
rect 1126 -1133 1230 -1128
rect 1082 -1183 1086 -1173
rect 1126 -1183 1131 -1133
rect 1257 -1137 1261 -1127
rect 1031 -1187 1045 -1183
rect 1039 -1188 1045 -1187
rect 1056 -1188 1074 -1183
rect 1082 -1188 1131 -1183
rect 1249 -1183 1253 -1177
rect 1274 -1183 1279 -1127
rect 1284 -1126 1287 -1122
rect 1291 -1126 1304 -1122
rect 1308 -1126 1311 -1122
rect 1284 -1128 1311 -1126
rect 1292 -1133 1296 -1128
rect 1300 -1183 1304 -1173
rect 1691 -1183 1696 -978
rect 1747 -979 1788 -974
rect 1796 -979 1904 -974
rect 1747 -982 1751 -979
rect 1796 -982 1800 -979
rect 1732 -986 1769 -982
rect 1732 -992 1736 -986
rect 1765 -992 1769 -986
rect 1899 -1000 1904 -979
rect 2134 -981 2161 -978
rect 2134 -985 2137 -981
rect 2141 -985 2154 -981
rect 2158 -985 2161 -981
rect 2134 -987 2161 -985
rect 2142 -992 2146 -987
rect 2031 -1000 2036 -998
rect 1788 -1008 1792 -1002
rect 1899 -1005 2036 -1000
rect 1780 -1009 1807 -1008
rect 1724 -1018 1728 -1012
rect 1757 -1018 1761 -1012
rect 1780 -1013 1781 -1009
rect 1785 -1013 1802 -1009
rect 1806 -1013 1807 -1009
rect 1780 -1014 1807 -1013
rect 1996 -1009 2002 -1008
rect 1996 -1013 1997 -1009
rect 2001 -1013 2002 -1009
rect 1996 -1016 2002 -1013
rect 2031 -1016 2036 -1005
rect 2091 -1011 2100 -1008
rect 2091 -1015 2093 -1011
rect 2097 -1015 2100 -1011
rect 2114 -1015 2127 -1012
rect 2091 -1016 2100 -1015
rect 1716 -1019 1743 -1018
rect 1716 -1023 1717 -1019
rect 1721 -1023 1738 -1019
rect 1742 -1023 1743 -1019
rect 1716 -1024 1743 -1023
rect 1749 -1019 1776 -1018
rect 1749 -1023 1750 -1019
rect 1754 -1023 1771 -1019
rect 1775 -1023 1776 -1019
rect 1749 -1024 1776 -1023
rect 1996 -1020 2008 -1016
rect 1996 -1030 2002 -1020
rect 2086 -1020 2100 -1016
rect 2028 -1028 2046 -1024
rect 2091 -1028 2100 -1020
rect 1996 -1034 1997 -1030
rect 2001 -1034 2002 -1030
rect 1996 -1035 2002 -1034
rect 2031 -1038 2036 -1028
rect 2091 -1032 2093 -1028
rect 2097 -1032 2100 -1028
rect 2091 -1035 2100 -1032
rect 2106 -1038 2110 -1035
rect 2060 -1042 2110 -1038
rect 1249 -1187 1263 -1183
rect 1257 -1188 1263 -1187
rect 1274 -1188 1292 -1183
rect 1300 -1188 1696 -1183
rect 1773 -1047 1779 -1046
rect 2060 -1047 2064 -1042
rect 1773 -1052 2064 -1047
rect 2114 -1048 2118 -1035
rect 2121 -1042 2127 -1015
rect 2150 -1042 2154 -1032
rect 2121 -1047 2142 -1042
rect 2150 -1047 2161 -1042
rect 995 -1199 1031 -1194
rect 1039 -1202 1043 -1188
rect 1082 -1191 1086 -1188
rect 229 -1213 233 -1203
rect 178 -1217 192 -1213
rect 186 -1218 192 -1217
rect 203 -1218 221 -1213
rect 229 -1218 335 -1213
rect 340 -1218 364 -1213
rect -3126 -1227 -3099 -1224
rect -3172 -1232 -3131 -1228
rect -3481 -1290 -3477 -1259
rect -3346 -1249 -3342 -1239
rect -3306 -1244 -3289 -1239
rect -3281 -1248 -3277 -1236
rect -3187 -1238 -3180 -1233
rect -3153 -1242 -3149 -1232
rect -3362 -1254 -3354 -1249
rect -3346 -1254 -3333 -1249
rect -3289 -1252 -3277 -1248
rect -3346 -1257 -3342 -1254
rect -3445 -1267 -3441 -1261
rect -3453 -1268 -3426 -1267
rect -3453 -1272 -3452 -1268
rect -3448 -1272 -3431 -1268
rect -3427 -1272 -3426 -1268
rect -3453 -1273 -3426 -1272
rect -3289 -1256 -3285 -1252
rect -3354 -1283 -3350 -1277
rect -3362 -1284 -3335 -1283
rect -3362 -1288 -3361 -1284
rect -3357 -1288 -3340 -1284
rect -3336 -1288 -3335 -1284
rect -3362 -1289 -3335 -1288
rect -3556 -1293 -3477 -1290
rect -3248 -1282 -3221 -1279
rect -3248 -1286 -3245 -1282
rect -3241 -1286 -3228 -1282
rect -3224 -1286 -3221 -1282
rect -3248 -1288 -3221 -1286
rect -3161 -1288 -3157 -1282
rect -3136 -1288 -3131 -1232
rect -3126 -1231 -3123 -1227
rect -3119 -1231 -3106 -1227
rect -3102 -1231 -3099 -1227
rect 57 -1229 178 -1224
rect -3126 -1233 -3099 -1231
rect 186 -1232 190 -1218
rect 229 -1221 233 -1218
rect -3118 -1238 -3114 -1233
rect 221 -1247 225 -1241
rect 1142 -1199 1249 -1194
rect 1074 -1217 1078 -1211
rect 1066 -1218 1093 -1217
rect 1066 -1222 1067 -1218
rect 1071 -1222 1088 -1218
rect 1092 -1222 1093 -1218
rect 1066 -1223 1093 -1222
rect 213 -1248 240 -1247
rect 1031 -1248 1035 -1242
rect 213 -1252 214 -1248
rect 218 -1252 235 -1248
rect 239 -1252 240 -1248
rect 213 -1253 240 -1252
rect 1023 -1249 1050 -1248
rect 1023 -1253 1024 -1249
rect 1028 -1253 1045 -1249
rect 1049 -1253 1050 -1249
rect 1023 -1254 1050 -1253
rect 1142 -1266 1147 -1199
rect 1257 -1202 1261 -1188
rect 1300 -1191 1304 -1188
rect 1292 -1217 1296 -1211
rect 1284 -1218 1311 -1217
rect 1284 -1222 1285 -1218
rect 1289 -1222 1306 -1218
rect 1310 -1222 1311 -1218
rect 1284 -1223 1311 -1222
rect 1249 -1248 1253 -1242
rect 1241 -1249 1268 -1248
rect 1241 -1253 1242 -1249
rect 1246 -1253 1263 -1249
rect 1267 -1253 1268 -1249
rect 1241 -1254 1268 -1253
rect 331 -1271 1147 -1266
rect 178 -1278 182 -1272
rect -3110 -1288 -3106 -1278
rect 170 -1279 197 -1278
rect 170 -1283 171 -1279
rect 175 -1283 192 -1279
rect 196 -1283 197 -1279
rect 170 -1284 197 -1283
rect 1773 -1288 1779 -1052
rect 1996 -1060 2002 -1059
rect 1996 -1064 1997 -1060
rect 2001 -1064 2002 -1060
rect 1996 -1067 2002 -1064
rect 2031 -1067 2036 -1052
rect 2091 -1062 2100 -1059
rect 2091 -1066 2093 -1062
rect 2097 -1066 2100 -1062
rect 2091 -1067 2100 -1066
rect 1996 -1071 2008 -1067
rect 1996 -1081 2002 -1071
rect 2086 -1071 2100 -1067
rect 2028 -1079 2046 -1075
rect 2091 -1079 2100 -1071
rect 1996 -1085 1997 -1081
rect 2001 -1085 2002 -1081
rect 1996 -1086 2002 -1085
rect 2031 -1099 2036 -1079
rect 2091 -1083 2093 -1079
rect 2097 -1083 2100 -1079
rect 2091 -1086 2100 -1083
rect 2150 -1050 2154 -1047
rect 2106 -1099 2110 -1068
rect 2142 -1076 2146 -1070
rect 2134 -1077 2161 -1076
rect 2134 -1081 2135 -1077
rect 2139 -1081 2156 -1077
rect 2160 -1081 2161 -1077
rect 2134 -1082 2161 -1081
rect 2031 -1102 2110 -1099
rect -3240 -1293 -3236 -1288
rect -3161 -1292 -3147 -1288
rect -3153 -1293 -3147 -1292
rect -3136 -1293 -3118 -1288
rect -3110 -1293 -3097 -1288
rect -3187 -1304 -3161 -1299
rect -3153 -1307 -3149 -1293
rect -3110 -1296 -3106 -1293
rect -3313 -1347 -3304 -1342
rect -3281 -1343 -3277 -1336
rect -3232 -1343 -3228 -1333
rect -3281 -1348 -3240 -1343
rect -3232 -1348 -3221 -1343
rect 344 -1294 1779 -1288
rect 344 -1299 350 -1294
rect 349 -1305 350 -1299
rect 344 -1313 350 -1305
rect 353 -1310 1212 -1305
rect 353 -1314 358 -1310
rect -3118 -1322 -3114 -1316
rect 353 -1322 358 -1319
rect -3126 -1323 -3099 -1322
rect -3126 -1327 -3125 -1323
rect -3121 -1327 -3104 -1323
rect -3100 -1327 -3099 -1323
rect -3126 -1328 -3099 -1327
rect 766 -1344 820 -1341
rect -3281 -1351 -3277 -1348
rect -3232 -1351 -3228 -1348
rect -3296 -1355 -3259 -1351
rect -3296 -1361 -3292 -1355
rect -3263 -1361 -3259 -1355
rect -3161 -1353 -3157 -1347
rect 766 -1348 769 -1344
rect 773 -1348 786 -1344
rect 790 -1348 796 -1344
rect 800 -1348 813 -1344
rect 817 -1348 820 -1344
rect 766 -1350 820 -1348
rect -3169 -1354 -3142 -1353
rect -3169 -1358 -3168 -1354
rect -3164 -1358 -3147 -1354
rect -3143 -1358 -3142 -1354
rect -3169 -1359 -3142 -1358
rect 774 -1355 778 -1350
rect 801 -1355 805 -1350
rect -3240 -1377 -3236 -1371
rect -3248 -1378 -3221 -1377
rect -3304 -1387 -3300 -1381
rect -3271 -1387 -3267 -1381
rect -3248 -1382 -3247 -1378
rect -3243 -1382 -3226 -1378
rect -3222 -1382 -3221 -1378
rect -3248 -1383 -3221 -1382
rect -3312 -1388 -3285 -1387
rect -3312 -1392 -3311 -1388
rect -3307 -1392 -3290 -1388
rect -3286 -1392 -3285 -1388
rect -3312 -1393 -3285 -1392
rect -3279 -1388 -3252 -1387
rect -3279 -1392 -3278 -1388
rect -3274 -1392 -3257 -1388
rect -3253 -1392 -3252 -1388
rect -3279 -1393 -3252 -1392
rect 782 -1415 786 -1395
rect 809 -1415 813 -1395
rect 828 -1414 855 -1411
rect 782 -1419 823 -1415
rect 349 -1425 774 -1420
rect 801 -1429 805 -1419
rect 793 -1475 797 -1469
rect 818 -1475 823 -1419
rect 828 -1418 831 -1414
rect 835 -1418 848 -1414
rect 852 -1418 855 -1414
rect 828 -1420 855 -1418
rect 836 -1425 840 -1420
rect 844 -1475 848 -1465
rect 793 -1479 807 -1475
rect 801 -1480 807 -1479
rect 818 -1480 836 -1475
rect 844 -1476 857 -1475
rect 844 -1480 1184 -1476
rect 340 -1491 793 -1486
rect 801 -1494 805 -1480
rect 844 -1483 848 -1480
rect 851 -1481 1184 -1480
rect 836 -1509 840 -1503
rect 828 -1510 855 -1509
rect 828 -1514 829 -1510
rect 833 -1514 850 -1510
rect 854 -1514 855 -1510
rect 828 -1515 855 -1514
rect 793 -1540 797 -1534
rect 785 -1541 812 -1540
rect 785 -1545 786 -1541
rect 790 -1545 807 -1541
rect 811 -1545 812 -1541
rect 785 -1546 812 -1545
rect 1003 -1574 1057 -1571
rect 1003 -1578 1006 -1574
rect 1010 -1578 1023 -1574
rect 1027 -1578 1033 -1574
rect 1037 -1578 1050 -1574
rect 1054 -1578 1057 -1574
rect 1003 -1580 1057 -1578
rect 1011 -1585 1015 -1580
rect 1038 -1585 1042 -1580
rect 243 -1598 270 -1595
rect 243 -1602 246 -1598
rect 250 -1602 263 -1598
rect 267 -1602 270 -1598
rect 243 -1604 270 -1602
rect 251 -1609 255 -1604
rect 140 -1617 145 -1615
rect -22 -1622 11 -1617
rect 16 -1622 145 -1617
rect 105 -1626 111 -1625
rect 105 -1630 106 -1626
rect 110 -1630 111 -1626
rect 105 -1633 111 -1630
rect 140 -1633 145 -1622
rect 200 -1628 209 -1625
rect 200 -1632 202 -1628
rect 206 -1632 209 -1628
rect 223 -1632 236 -1629
rect 200 -1633 209 -1632
rect 105 -1637 117 -1633
rect 105 -1647 111 -1637
rect 195 -1637 209 -1633
rect 137 -1645 155 -1641
rect 200 -1645 209 -1637
rect 105 -1651 106 -1647
rect 110 -1651 111 -1647
rect 105 -1652 111 -1651
rect 140 -1655 145 -1645
rect 200 -1649 202 -1645
rect 206 -1649 209 -1645
rect 200 -1652 209 -1649
rect 215 -1655 219 -1652
rect 169 -1659 219 -1655
rect 169 -1664 173 -1659
rect -19 -1669 173 -1664
rect 223 -1665 227 -1652
rect 230 -1659 236 -1632
rect 767 -1627 821 -1624
rect 767 -1631 770 -1627
rect 774 -1631 787 -1627
rect 791 -1631 797 -1627
rect 801 -1631 814 -1627
rect 818 -1631 821 -1627
rect 767 -1633 821 -1631
rect 259 -1659 263 -1649
rect 775 -1638 779 -1633
rect 802 -1638 806 -1633
rect 230 -1664 251 -1659
rect 259 -1664 344 -1659
rect 349 -1664 378 -1659
rect 66 -1884 71 -1669
rect 105 -1677 111 -1676
rect 105 -1681 106 -1677
rect 110 -1681 111 -1677
rect 105 -1684 111 -1681
rect 140 -1684 145 -1669
rect 200 -1679 209 -1676
rect 200 -1683 202 -1679
rect 206 -1683 209 -1679
rect 200 -1684 209 -1683
rect 105 -1688 117 -1684
rect 105 -1698 111 -1688
rect 195 -1688 209 -1684
rect 137 -1696 155 -1692
rect 200 -1696 209 -1688
rect 105 -1702 106 -1698
rect 110 -1702 111 -1698
rect 105 -1703 111 -1702
rect 140 -1716 145 -1696
rect 200 -1700 202 -1696
rect 206 -1700 209 -1696
rect 200 -1703 209 -1700
rect 259 -1667 263 -1664
rect 215 -1716 219 -1685
rect 1019 -1645 1023 -1625
rect 1046 -1645 1050 -1625
rect 1065 -1644 1092 -1641
rect 1019 -1649 1060 -1645
rect 1004 -1651 1011 -1650
rect 251 -1693 255 -1687
rect 243 -1694 270 -1693
rect 243 -1698 244 -1694
rect 248 -1698 265 -1694
rect 269 -1698 270 -1694
rect 243 -1699 270 -1698
rect 783 -1698 787 -1678
rect 810 -1698 814 -1678
rect 943 -1655 1011 -1651
rect 943 -1656 1009 -1655
rect 829 -1697 856 -1694
rect 783 -1702 824 -1698
rect 349 -1708 775 -1703
rect 802 -1712 806 -1702
rect 140 -1719 219 -1716
rect 160 -1742 214 -1739
rect 160 -1746 163 -1742
rect 167 -1746 180 -1742
rect 184 -1746 190 -1742
rect 194 -1746 207 -1742
rect 211 -1746 214 -1742
rect 160 -1748 214 -1746
rect 168 -1753 172 -1748
rect 195 -1753 199 -1748
rect 794 -1758 798 -1752
rect 819 -1758 824 -1702
rect 829 -1701 832 -1697
rect 836 -1701 849 -1697
rect 853 -1701 856 -1697
rect 829 -1703 856 -1701
rect 837 -1708 841 -1703
rect 845 -1758 849 -1748
rect 943 -1758 948 -1656
rect 1038 -1659 1042 -1649
rect 1030 -1705 1034 -1699
rect 1055 -1705 1060 -1649
rect 1065 -1648 1068 -1644
rect 1072 -1648 1085 -1644
rect 1089 -1648 1092 -1644
rect 1065 -1650 1092 -1648
rect 1073 -1655 1077 -1650
rect 1179 -1668 1184 -1481
rect 1207 -1565 1212 -1310
rect 1417 -1471 1444 -1468
rect 1417 -1475 1420 -1471
rect 1424 -1475 1437 -1471
rect 1441 -1475 1444 -1471
rect 1417 -1477 1444 -1475
rect 1425 -1482 1429 -1477
rect 1207 -1570 1425 -1565
rect 1433 -1574 1437 -1562
rect 1425 -1578 1437 -1574
rect 1425 -1582 1429 -1578
rect 1466 -1608 1493 -1605
rect 1466 -1612 1469 -1608
rect 1473 -1612 1486 -1608
rect 1490 -1612 1493 -1608
rect 1466 -1614 1493 -1612
rect 1474 -1619 1478 -1614
rect 1714 -1624 1741 -1621
rect 1714 -1628 1717 -1624
rect 1721 -1628 1734 -1624
rect 1738 -1628 1741 -1624
rect 1714 -1630 1741 -1628
rect 1179 -1673 1410 -1668
rect 1433 -1669 1437 -1662
rect 1482 -1669 1486 -1659
rect 1722 -1635 1726 -1630
rect 1433 -1674 1474 -1669
rect 1482 -1674 1710 -1669
rect 1433 -1677 1437 -1674
rect 1482 -1677 1486 -1674
rect 1418 -1681 1455 -1677
rect 1418 -1687 1422 -1681
rect 1451 -1687 1455 -1681
rect 1081 -1705 1085 -1695
rect 1030 -1709 1044 -1705
rect 1038 -1710 1044 -1709
rect 1055 -1710 1073 -1705
rect 1081 -1706 1094 -1705
rect 1081 -1710 1175 -1706
rect 794 -1762 808 -1758
rect 802 -1763 808 -1762
rect 819 -1763 837 -1758
rect 845 -1763 948 -1758
rect 964 -1721 1030 -1716
rect 331 -1774 794 -1769
rect 802 -1777 806 -1763
rect 845 -1766 849 -1763
rect 176 -1813 180 -1793
rect 203 -1813 207 -1793
rect 222 -1812 249 -1809
rect 176 -1817 217 -1813
rect 104 -1823 168 -1818
rect 195 -1827 199 -1817
rect 187 -1873 191 -1867
rect 212 -1873 217 -1817
rect 222 -1816 225 -1812
rect 229 -1816 242 -1812
rect 246 -1816 249 -1812
rect 222 -1818 249 -1816
rect 837 -1792 841 -1786
rect 829 -1793 856 -1792
rect 829 -1797 830 -1793
rect 834 -1797 851 -1793
rect 855 -1797 856 -1793
rect 829 -1798 856 -1797
rect 230 -1823 234 -1818
rect 794 -1823 798 -1817
rect 786 -1824 813 -1823
rect 786 -1828 787 -1824
rect 791 -1828 808 -1824
rect 812 -1828 813 -1824
rect 786 -1829 813 -1828
rect 964 -1840 969 -1721
rect 1038 -1724 1042 -1710
rect 1081 -1713 1085 -1710
rect 1088 -1711 1175 -1710
rect 1073 -1739 1077 -1733
rect 1065 -1740 1092 -1739
rect 1065 -1744 1066 -1740
rect 1070 -1744 1087 -1740
rect 1091 -1744 1092 -1740
rect 1065 -1745 1092 -1744
rect 1030 -1770 1034 -1764
rect 1022 -1771 1049 -1770
rect 1022 -1775 1023 -1771
rect 1027 -1775 1044 -1771
rect 1048 -1775 1049 -1771
rect 1022 -1776 1049 -1775
rect 1012 -1785 1066 -1782
rect 1012 -1789 1015 -1785
rect 1019 -1789 1032 -1785
rect 1036 -1789 1042 -1785
rect 1046 -1789 1059 -1785
rect 1063 -1789 1066 -1785
rect 1012 -1791 1066 -1789
rect 1020 -1796 1024 -1791
rect 1047 -1796 1051 -1791
rect 322 -1845 969 -1840
rect 1028 -1856 1032 -1836
rect 1055 -1856 1059 -1836
rect 1074 -1855 1101 -1852
rect 1028 -1860 1069 -1856
rect 1013 -1862 1020 -1861
rect 238 -1873 242 -1863
rect 949 -1866 1020 -1862
rect 949 -1867 1016 -1866
rect 187 -1877 201 -1873
rect 195 -1878 201 -1877
rect 212 -1878 230 -1873
rect 238 -1878 353 -1873
rect 358 -1878 391 -1873
rect 66 -1889 187 -1884
rect 195 -1892 199 -1878
rect 238 -1881 242 -1878
rect 763 -1898 817 -1895
rect 230 -1907 234 -1901
rect 763 -1902 766 -1898
rect 770 -1902 783 -1898
rect 787 -1902 793 -1898
rect 797 -1902 810 -1898
rect 814 -1902 817 -1898
rect 763 -1904 817 -1902
rect 222 -1908 249 -1907
rect 222 -1912 223 -1908
rect 227 -1912 244 -1908
rect 248 -1912 249 -1908
rect 222 -1913 249 -1912
rect 771 -1909 775 -1904
rect 798 -1909 802 -1904
rect 187 -1938 191 -1932
rect 179 -1939 206 -1938
rect 179 -1943 180 -1939
rect 184 -1943 201 -1939
rect 205 -1943 206 -1939
rect 179 -1944 206 -1943
rect 779 -1969 783 -1949
rect 806 -1969 810 -1949
rect 825 -1968 852 -1965
rect 779 -1973 820 -1969
rect 304 -1979 771 -1974
rect 798 -1983 802 -1973
rect 790 -2029 794 -2023
rect 815 -2029 820 -1973
rect 825 -1972 828 -1968
rect 832 -1972 845 -1968
rect 849 -1972 852 -1968
rect 825 -1974 852 -1972
rect 833 -1979 837 -1974
rect 841 -2029 845 -2019
rect 949 -2029 954 -1867
rect 1047 -1870 1051 -1860
rect 1039 -1916 1043 -1910
rect 1064 -1916 1069 -1860
rect 1074 -1859 1077 -1855
rect 1081 -1859 1094 -1855
rect 1098 -1859 1101 -1855
rect 1074 -1861 1101 -1859
rect 1082 -1866 1086 -1861
rect 1170 -1865 1175 -1711
rect 1474 -1703 1478 -1697
rect 1466 -1704 1493 -1703
rect 1410 -1713 1414 -1707
rect 1443 -1713 1447 -1707
rect 1466 -1708 1467 -1704
rect 1471 -1708 1488 -1704
rect 1492 -1708 1493 -1704
rect 1466 -1709 1493 -1708
rect 1402 -1714 1429 -1713
rect 1402 -1718 1403 -1714
rect 1407 -1718 1424 -1714
rect 1428 -1718 1429 -1714
rect 1402 -1719 1429 -1718
rect 1435 -1714 1462 -1713
rect 1435 -1718 1436 -1714
rect 1440 -1718 1457 -1714
rect 1461 -1718 1462 -1714
rect 1435 -1719 1462 -1718
rect 1705 -1718 1710 -1674
rect 2132 -1689 2159 -1686
rect 2132 -1693 2135 -1689
rect 2139 -1693 2152 -1689
rect 2156 -1693 2159 -1689
rect 2132 -1695 2159 -1693
rect 2140 -1700 2144 -1695
rect 1705 -1723 1722 -1718
rect 1730 -1727 1734 -1715
rect 1722 -1731 1734 -1727
rect 1899 -1708 1999 -1705
rect 2029 -1708 2034 -1706
rect 1899 -1710 2034 -1708
rect 1722 -1735 1726 -1731
rect 1428 -1771 1455 -1768
rect 1428 -1775 1431 -1771
rect 1435 -1775 1448 -1771
rect 1452 -1775 1455 -1771
rect 1428 -1777 1455 -1775
rect 1436 -1782 1440 -1777
rect 1763 -1761 1790 -1758
rect 1763 -1765 1766 -1761
rect 1770 -1765 1783 -1761
rect 1787 -1765 1790 -1761
rect 1763 -1767 1790 -1765
rect 1771 -1772 1775 -1767
rect 1170 -1870 1436 -1865
rect 1444 -1874 1448 -1862
rect 1090 -1916 1094 -1906
rect 1436 -1878 1448 -1874
rect 1679 -1826 1707 -1821
rect 1730 -1822 1734 -1815
rect 1779 -1822 1783 -1812
rect 1899 -1822 1904 -1710
rect 1994 -1713 2034 -1710
rect 1994 -1717 2000 -1716
rect 1994 -1721 1995 -1717
rect 1999 -1721 2000 -1717
rect 1994 -1724 2000 -1721
rect 2029 -1724 2034 -1713
rect 2089 -1719 2098 -1716
rect 2089 -1723 2091 -1719
rect 2095 -1723 2098 -1719
rect 2112 -1723 2125 -1720
rect 2089 -1724 2098 -1723
rect 1994 -1728 2006 -1724
rect 1994 -1738 2000 -1728
rect 2084 -1728 2098 -1724
rect 2026 -1736 2044 -1732
rect 2089 -1736 2098 -1728
rect 1994 -1742 1995 -1738
rect 1999 -1742 2000 -1738
rect 1994 -1743 2000 -1742
rect 2029 -1746 2034 -1736
rect 2089 -1740 2091 -1736
rect 2095 -1740 2098 -1736
rect 2089 -1743 2098 -1740
rect 2104 -1746 2108 -1743
rect 2058 -1750 2108 -1746
rect 2058 -1755 2062 -1750
rect 1436 -1882 1440 -1878
rect 1039 -1920 1053 -1916
rect 1047 -1921 1053 -1920
rect 1064 -1921 1082 -1916
rect 1090 -1921 1128 -1916
rect 1013 -1928 1039 -1927
rect 790 -2033 804 -2029
rect 798 -2034 804 -2033
rect 815 -2034 833 -2029
rect 841 -2034 954 -2029
rect 988 -1932 1039 -1928
rect 988 -1933 1029 -1932
rect 307 -2045 308 -2040
rect 313 -2045 790 -2040
rect 798 -2048 802 -2034
rect 841 -2037 845 -2034
rect 833 -2063 837 -2057
rect 825 -2064 852 -2063
rect 825 -2068 826 -2064
rect 830 -2068 847 -2064
rect 851 -2068 852 -2064
rect 825 -2069 852 -2068
rect 790 -2094 794 -2088
rect 782 -2095 809 -2094
rect 782 -2099 783 -2095
rect 787 -2099 804 -2095
rect 808 -2099 809 -2095
rect 782 -2100 809 -2099
rect 751 -2147 805 -2144
rect 751 -2151 754 -2147
rect 758 -2151 771 -2147
rect 775 -2151 781 -2147
rect 785 -2151 798 -2147
rect 802 -2151 805 -2147
rect 751 -2153 805 -2151
rect 759 -2158 763 -2153
rect 786 -2158 790 -2153
rect 767 -2218 771 -2198
rect 794 -2218 798 -2198
rect 813 -2217 840 -2214
rect 767 -2222 808 -2218
rect 343 -2228 344 -2223
rect 349 -2228 759 -2223
rect 786 -2232 790 -2222
rect 778 -2278 782 -2272
rect 803 -2278 808 -2222
rect 813 -2221 816 -2217
rect 820 -2221 833 -2217
rect 837 -2221 840 -2217
rect 813 -2223 840 -2221
rect 821 -2228 825 -2223
rect 829 -2278 833 -2268
rect 988 -2278 993 -1933
rect 1047 -1935 1051 -1921
rect 1090 -1924 1094 -1921
rect 1082 -1950 1086 -1944
rect 1074 -1951 1101 -1950
rect 1074 -1955 1075 -1951
rect 1079 -1955 1096 -1951
rect 1100 -1955 1101 -1951
rect 1074 -1956 1101 -1955
rect 1123 -1968 1128 -1921
rect 1477 -1908 1504 -1905
rect 1477 -1912 1480 -1908
rect 1484 -1912 1497 -1908
rect 1501 -1912 1504 -1908
rect 1477 -1914 1504 -1912
rect 1485 -1919 1489 -1914
rect 1123 -1973 1421 -1968
rect 1444 -1969 1448 -1962
rect 1493 -1969 1497 -1959
rect 1679 -1969 1684 -1826
rect 1730 -1827 1771 -1822
rect 1779 -1827 1904 -1822
rect 1908 -1760 2062 -1755
rect 2112 -1756 2116 -1743
rect 2119 -1750 2125 -1723
rect 2148 -1750 2152 -1740
rect 2119 -1755 2140 -1750
rect 2148 -1755 2159 -1750
rect 1730 -1830 1734 -1827
rect 1779 -1830 1783 -1827
rect 1715 -1834 1752 -1830
rect 1715 -1840 1719 -1834
rect 1748 -1840 1752 -1834
rect 1771 -1856 1775 -1850
rect 1763 -1857 1790 -1856
rect 1707 -1866 1711 -1860
rect 1740 -1866 1744 -1860
rect 1763 -1861 1764 -1857
rect 1768 -1861 1785 -1857
rect 1789 -1861 1790 -1857
rect 1763 -1862 1790 -1861
rect 1699 -1867 1726 -1866
rect 1699 -1871 1700 -1867
rect 1704 -1871 1721 -1867
rect 1725 -1871 1726 -1867
rect 1699 -1872 1726 -1871
rect 1732 -1867 1759 -1866
rect 1732 -1871 1733 -1867
rect 1737 -1871 1754 -1867
rect 1758 -1871 1759 -1867
rect 1732 -1872 1759 -1871
rect 1444 -1974 1485 -1969
rect 1493 -1974 1684 -1969
rect 1039 -1981 1043 -1975
rect 1444 -1977 1448 -1974
rect 1493 -1977 1497 -1974
rect 1429 -1981 1466 -1977
rect 1031 -1982 1058 -1981
rect 1031 -1986 1032 -1982
rect 1036 -1986 1053 -1982
rect 1057 -1986 1058 -1982
rect 1031 -1987 1058 -1986
rect 1429 -1987 1433 -1981
rect 1462 -1987 1466 -1981
rect 1485 -2003 1489 -1997
rect 1477 -2004 1504 -2003
rect 1421 -2013 1425 -2007
rect 1454 -2013 1458 -2007
rect 1477 -2008 1478 -2004
rect 1482 -2008 1499 -2004
rect 1503 -2008 1504 -2004
rect 1477 -2009 1504 -2008
rect 1413 -2014 1440 -2013
rect 1413 -2018 1414 -2014
rect 1418 -2018 1435 -2014
rect 1439 -2018 1440 -2014
rect 1413 -2019 1440 -2018
rect 1446 -2014 1473 -2013
rect 1446 -2018 1447 -2014
rect 1451 -2018 1468 -2014
rect 1472 -2018 1473 -2014
rect 1446 -2019 1473 -2018
rect 1908 -2098 1913 -1760
rect 1994 -1768 2000 -1767
rect 1994 -1772 1995 -1768
rect 1999 -1772 2000 -1768
rect 1994 -1775 2000 -1772
rect 2029 -1775 2034 -1760
rect 2089 -1770 2098 -1767
rect 2089 -1774 2091 -1770
rect 2095 -1774 2098 -1770
rect 2089 -1775 2098 -1774
rect 1994 -1779 2006 -1775
rect 1994 -1789 2000 -1779
rect 2084 -1779 2098 -1775
rect 2026 -1787 2044 -1783
rect 2089 -1787 2098 -1779
rect 1994 -1793 1995 -1789
rect 1999 -1793 2000 -1789
rect 1994 -1794 2000 -1793
rect 2029 -1807 2034 -1787
rect 2089 -1791 2091 -1787
rect 2095 -1791 2098 -1787
rect 2089 -1794 2098 -1791
rect 2148 -1758 2152 -1755
rect 2104 -1807 2108 -1776
rect 2140 -1784 2144 -1778
rect 2132 -1785 2159 -1784
rect 2132 -1789 2133 -1785
rect 2137 -1789 2154 -1785
rect 2158 -1789 2159 -1785
rect 2132 -1790 2159 -1789
rect 2029 -1810 2108 -1807
rect 778 -2282 792 -2278
rect 786 -2283 792 -2282
rect 803 -2283 821 -2278
rect 829 -2283 993 -2278
rect 1016 -2103 1913 -2098
rect 331 -2294 778 -2289
rect 786 -2297 790 -2283
rect 829 -2286 833 -2283
rect 821 -2312 825 -2306
rect 813 -2313 840 -2312
rect 813 -2317 814 -2313
rect 818 -2317 835 -2313
rect 839 -2317 840 -2313
rect 813 -2318 840 -2317
rect 778 -2343 782 -2337
rect 770 -2344 797 -2343
rect 770 -2348 771 -2344
rect 775 -2348 792 -2344
rect 796 -2348 797 -2344
rect 770 -2349 797 -2348
rect 1016 -2378 1021 -2103
rect 360 -2383 362 -2378
rect 367 -2383 1021 -2378
rect 523 -2460 1409 -2455
rect 240 -2473 267 -2470
rect 240 -2477 243 -2473
rect 247 -2477 260 -2473
rect 264 -2477 267 -2473
rect 240 -2479 267 -2477
rect 248 -2484 252 -2479
rect 137 -2492 142 -2490
rect -25 -2497 8 -2492
rect 13 -2497 142 -2492
rect 102 -2501 108 -2500
rect 102 -2505 103 -2501
rect 107 -2505 108 -2501
rect 102 -2508 108 -2505
rect 137 -2508 142 -2497
rect 197 -2503 206 -2500
rect 197 -2507 199 -2503
rect 203 -2507 206 -2503
rect 220 -2507 233 -2504
rect 197 -2508 206 -2507
rect 102 -2512 114 -2508
rect 102 -2522 108 -2512
rect 192 -2512 206 -2508
rect 134 -2520 152 -2516
rect 197 -2520 206 -2512
rect 102 -2526 103 -2522
rect 107 -2526 108 -2522
rect 102 -2527 108 -2526
rect 137 -2530 142 -2520
rect 197 -2524 199 -2520
rect 203 -2524 206 -2520
rect 197 -2527 206 -2524
rect 212 -2530 216 -2527
rect 166 -2534 216 -2530
rect 166 -2539 170 -2534
rect -22 -2544 170 -2539
rect 220 -2540 224 -2527
rect 227 -2534 233 -2507
rect 256 -2534 260 -2524
rect 227 -2539 248 -2534
rect 256 -2539 362 -2534
rect 367 -2539 387 -2534
rect 63 -2759 68 -2544
rect 102 -2552 108 -2551
rect 102 -2556 103 -2552
rect 107 -2556 108 -2552
rect 102 -2559 108 -2556
rect 137 -2559 142 -2544
rect 197 -2554 206 -2551
rect 197 -2558 199 -2554
rect 203 -2558 206 -2554
rect 197 -2559 206 -2558
rect 102 -2563 114 -2559
rect 102 -2573 108 -2563
rect 192 -2563 206 -2559
rect 134 -2571 152 -2567
rect 197 -2571 206 -2563
rect 102 -2577 103 -2573
rect 107 -2577 108 -2573
rect 102 -2578 108 -2577
rect 137 -2591 142 -2571
rect 197 -2575 199 -2571
rect 203 -2575 206 -2571
rect 197 -2578 206 -2575
rect 256 -2542 260 -2539
rect 212 -2591 216 -2560
rect 248 -2568 252 -2562
rect 240 -2569 267 -2568
rect 240 -2573 241 -2569
rect 245 -2573 262 -2569
rect 266 -2573 267 -2569
rect 240 -2574 267 -2573
rect 137 -2594 216 -2591
rect 157 -2617 211 -2614
rect 157 -2621 160 -2617
rect 164 -2621 177 -2617
rect 181 -2621 187 -2617
rect 191 -2621 204 -2617
rect 208 -2621 211 -2617
rect 157 -2623 211 -2621
rect 165 -2628 169 -2623
rect 192 -2628 196 -2623
rect 173 -2688 177 -2668
rect 200 -2688 204 -2668
rect 219 -2687 246 -2684
rect 173 -2692 214 -2688
rect 101 -2698 165 -2693
rect 192 -2702 196 -2692
rect 184 -2748 188 -2742
rect 209 -2748 214 -2692
rect 219 -2691 222 -2687
rect 226 -2691 239 -2687
rect 243 -2691 246 -2687
rect 219 -2693 246 -2691
rect 227 -2698 231 -2693
rect 235 -2748 239 -2738
rect 523 -2748 528 -2460
rect 1011 -2491 1379 -2486
rect 792 -2496 846 -2493
rect 792 -2500 795 -2496
rect 799 -2500 812 -2496
rect 816 -2500 822 -2496
rect 826 -2500 839 -2496
rect 843 -2500 846 -2496
rect 792 -2502 846 -2500
rect 800 -2507 804 -2502
rect 827 -2507 831 -2502
rect 808 -2567 812 -2547
rect 835 -2567 839 -2547
rect 854 -2566 881 -2563
rect 808 -2571 849 -2567
rect 184 -2752 198 -2748
rect 192 -2753 198 -2752
rect 209 -2753 227 -2748
rect 235 -2753 528 -2748
rect 537 -2577 800 -2572
rect 63 -2764 184 -2759
rect 192 -2767 196 -2753
rect 235 -2756 239 -2753
rect 537 -2765 542 -2577
rect 827 -2581 831 -2571
rect 819 -2627 823 -2621
rect 844 -2627 849 -2571
rect 854 -2570 857 -2566
rect 861 -2570 874 -2566
rect 878 -2570 881 -2566
rect 854 -2572 881 -2570
rect 862 -2577 866 -2572
rect 870 -2627 874 -2617
rect 1011 -2627 1016 -2491
rect 1127 -2548 1181 -2545
rect 1127 -2552 1130 -2548
rect 1134 -2552 1147 -2548
rect 1151 -2552 1157 -2548
rect 1161 -2552 1174 -2548
rect 1178 -2552 1181 -2548
rect 1127 -2554 1181 -2552
rect 1135 -2559 1139 -2554
rect 1162 -2559 1166 -2554
rect 1143 -2619 1147 -2599
rect 1170 -2619 1174 -2599
rect 1189 -2618 1216 -2615
rect 1143 -2623 1184 -2619
rect 819 -2631 833 -2627
rect 827 -2632 833 -2631
rect 844 -2632 862 -2627
rect 870 -2632 1016 -2627
rect 1124 -2629 1135 -2624
rect 352 -2770 353 -2765
rect 358 -2770 542 -2765
rect 550 -2643 819 -2638
rect 550 -2774 555 -2643
rect 827 -2646 831 -2632
rect 870 -2635 874 -2632
rect 1124 -2642 1132 -2629
rect 1162 -2633 1166 -2623
rect 1063 -2644 1132 -2642
rect 1016 -2649 1132 -2644
rect 862 -2661 866 -2655
rect 854 -2662 881 -2661
rect 854 -2666 855 -2662
rect 859 -2666 876 -2662
rect 880 -2666 881 -2662
rect 854 -2667 881 -2666
rect 819 -2692 823 -2686
rect 811 -2693 838 -2692
rect 811 -2697 812 -2693
rect 816 -2697 833 -2693
rect 837 -2697 838 -2693
rect 811 -2698 838 -2697
rect 227 -2782 231 -2776
rect 367 -2779 555 -2774
rect 793 -2779 847 -2776
rect 219 -2783 246 -2782
rect 219 -2787 220 -2783
rect 224 -2787 241 -2783
rect 245 -2787 246 -2783
rect 793 -2783 796 -2779
rect 800 -2783 813 -2779
rect 817 -2783 823 -2779
rect 827 -2783 840 -2779
rect 844 -2783 847 -2779
rect 793 -2785 847 -2783
rect 219 -2788 246 -2787
rect 801 -2790 805 -2785
rect 828 -2790 832 -2785
rect 184 -2813 188 -2807
rect 176 -2814 203 -2813
rect 176 -2818 177 -2814
rect 181 -2818 198 -2814
rect 202 -2818 203 -2814
rect 176 -2819 203 -2818
rect 809 -2850 813 -2830
rect 836 -2850 840 -2830
rect 855 -2849 882 -2846
rect 809 -2854 850 -2850
rect 361 -2860 362 -2855
rect 367 -2860 801 -2855
rect 828 -2864 832 -2854
rect 820 -2910 824 -2904
rect 845 -2910 850 -2854
rect 855 -2853 858 -2849
rect 862 -2853 875 -2849
rect 879 -2853 882 -2849
rect 855 -2855 882 -2853
rect 863 -2860 867 -2855
rect 871 -2910 875 -2900
rect 1016 -2910 1021 -2649
rect 1063 -2650 1132 -2649
rect 1154 -2679 1158 -2673
rect 1179 -2679 1184 -2623
rect 1189 -2622 1192 -2618
rect 1196 -2622 1209 -2618
rect 1213 -2622 1216 -2618
rect 1189 -2624 1216 -2622
rect 1197 -2629 1201 -2624
rect 1205 -2679 1209 -2669
rect 1154 -2683 1168 -2679
rect 1162 -2684 1168 -2683
rect 1179 -2684 1197 -2679
rect 1205 -2684 1363 -2679
rect 820 -2914 834 -2910
rect 828 -2915 834 -2914
rect 845 -2915 863 -2910
rect 871 -2915 1021 -2910
rect 1053 -2695 1154 -2690
rect 343 -2926 344 -2921
rect 349 -2926 820 -2921
rect 828 -2929 832 -2915
rect 871 -2918 875 -2915
rect 863 -2944 867 -2938
rect 855 -2945 882 -2944
rect 855 -2949 856 -2945
rect 860 -2949 877 -2945
rect 881 -2949 882 -2945
rect 855 -2950 882 -2949
rect 820 -2975 824 -2969
rect 812 -2976 839 -2975
rect 812 -2980 813 -2976
rect 817 -2980 834 -2976
rect 838 -2980 839 -2976
rect 812 -2981 839 -2980
rect 1053 -2995 1058 -2695
rect 1162 -2698 1166 -2684
rect 1205 -2687 1209 -2684
rect 1197 -2713 1201 -2707
rect 1189 -2714 1216 -2713
rect 1189 -2718 1190 -2714
rect 1194 -2718 1211 -2714
rect 1215 -2718 1216 -2714
rect 1189 -2719 1216 -2718
rect 1154 -2744 1158 -2738
rect 1146 -2745 1173 -2744
rect 1146 -2749 1147 -2745
rect 1151 -2749 1168 -2745
rect 1172 -2749 1173 -2745
rect 1146 -2750 1173 -2749
rect 1128 -2831 1182 -2828
rect 1128 -2835 1131 -2831
rect 1135 -2835 1148 -2831
rect 1152 -2835 1158 -2831
rect 1162 -2835 1175 -2831
rect 1179 -2835 1182 -2831
rect 1128 -2837 1182 -2835
rect 1136 -2842 1140 -2837
rect 1163 -2842 1167 -2837
rect 1144 -2902 1148 -2882
rect 1171 -2902 1175 -2882
rect 1190 -2901 1217 -2898
rect 1144 -2906 1185 -2902
rect 334 -3000 335 -2995
rect 340 -3000 1058 -2995
rect 1064 -2912 1136 -2907
rect 1064 -3013 1069 -2912
rect 1163 -2916 1167 -2906
rect 1155 -2962 1159 -2956
rect 1180 -2962 1185 -2906
rect 1190 -2905 1193 -2901
rect 1197 -2905 1210 -2901
rect 1214 -2905 1217 -2901
rect 1190 -2907 1217 -2905
rect 1198 -2912 1202 -2907
rect 1206 -2962 1210 -2952
rect 1155 -2966 1169 -2962
rect 1163 -2967 1169 -2966
rect 1180 -2967 1198 -2962
rect 1206 -2967 1346 -2962
rect 897 -3018 1069 -3013
rect 1081 -2978 1155 -2973
rect 789 -3050 843 -3047
rect 789 -3054 792 -3050
rect 796 -3054 809 -3050
rect 813 -3054 819 -3050
rect 823 -3054 836 -3050
rect 840 -3054 843 -3050
rect 789 -3056 843 -3054
rect 797 -3061 801 -3056
rect 824 -3061 828 -3056
rect 805 -3121 809 -3101
rect 832 -3121 836 -3101
rect 851 -3120 878 -3117
rect 805 -3125 846 -3121
rect 367 -3131 797 -3126
rect 824 -3135 828 -3125
rect 816 -3181 820 -3175
rect 841 -3181 846 -3125
rect 851 -3124 854 -3120
rect 858 -3124 871 -3120
rect 875 -3124 878 -3120
rect 851 -3126 878 -3124
rect 859 -3131 863 -3126
rect 867 -3181 871 -3171
rect 897 -3181 902 -3018
rect 1081 -3035 1086 -2978
rect 1163 -2981 1167 -2967
rect 1206 -2970 1210 -2967
rect 1198 -2996 1202 -2990
rect 1190 -2997 1217 -2996
rect 1190 -3001 1191 -2997
rect 1195 -3001 1212 -2997
rect 1216 -3001 1217 -2997
rect 1190 -3002 1217 -3001
rect 1155 -3027 1159 -3021
rect 1147 -3028 1174 -3027
rect 1147 -3032 1148 -3028
rect 1152 -3032 1169 -3028
rect 1173 -3032 1174 -3028
rect 1147 -3033 1174 -3032
rect 816 -3185 830 -3181
rect 824 -3186 830 -3185
rect 841 -3186 859 -3181
rect 867 -3186 902 -3181
rect 911 -3040 1086 -3035
rect 343 -3197 344 -3192
rect 349 -3197 816 -3192
rect 824 -3200 828 -3186
rect 867 -3189 871 -3186
rect 859 -3215 863 -3209
rect 851 -3216 878 -3215
rect 851 -3220 852 -3216
rect 856 -3220 873 -3216
rect 877 -3220 878 -3216
rect 851 -3221 878 -3220
rect 816 -3246 820 -3240
rect 808 -3247 835 -3246
rect 808 -3251 809 -3247
rect 813 -3251 830 -3247
rect 834 -3251 835 -3247
rect 808 -3252 835 -3251
rect 777 -3299 831 -3296
rect 777 -3303 780 -3299
rect 784 -3303 797 -3299
rect 801 -3303 807 -3299
rect 811 -3303 824 -3299
rect 828 -3303 831 -3299
rect 777 -3305 831 -3303
rect 785 -3310 789 -3305
rect 812 -3310 816 -3305
rect 793 -3370 797 -3350
rect 820 -3370 824 -3350
rect 839 -3369 866 -3366
rect 793 -3374 834 -3370
rect 322 -3380 785 -3375
rect 812 -3384 816 -3374
rect 804 -3430 808 -3424
rect 829 -3430 834 -3374
rect 839 -3373 842 -3369
rect 846 -3373 859 -3369
rect 863 -3373 866 -3369
rect 839 -3375 866 -3373
rect 847 -3380 851 -3375
rect 855 -3430 859 -3420
rect 911 -3430 916 -3040
rect 1341 -3075 1346 -2967
rect 1358 -2972 1363 -2684
rect 1374 -2686 1379 -2491
rect 1404 -2583 1409 -2460
rect 1457 -2489 1484 -2486
rect 1457 -2493 1460 -2489
rect 1464 -2493 1477 -2489
rect 1481 -2493 1484 -2489
rect 1457 -2495 1484 -2493
rect 1465 -2500 1469 -2495
rect 2192 -2513 2219 -2510
rect 2192 -2517 2195 -2513
rect 2199 -2517 2212 -2513
rect 2216 -2517 2219 -2513
rect 2192 -2519 2219 -2517
rect 1404 -2588 1465 -2583
rect 1404 -2589 1409 -2588
rect 1473 -2592 1477 -2580
rect 1465 -2596 1477 -2592
rect 2200 -2524 2204 -2519
rect 1465 -2600 1469 -2596
rect 2183 -2608 2200 -2607
rect 2021 -2612 2200 -2608
rect 2021 -2613 2185 -2612
rect 1506 -2626 1533 -2623
rect 1506 -2630 1509 -2626
rect 1513 -2630 1526 -2626
rect 1530 -2630 1533 -2626
rect 1506 -2632 1533 -2630
rect 1514 -2637 1518 -2632
rect 1374 -2691 1450 -2686
rect 1473 -2687 1477 -2680
rect 1522 -2687 1526 -2677
rect 2021 -2687 2026 -2613
rect 2208 -2616 2212 -2604
rect 1473 -2692 1514 -2687
rect 1522 -2692 2026 -2687
rect 2200 -2620 2212 -2616
rect 2200 -2624 2204 -2620
rect 1473 -2695 1477 -2692
rect 1522 -2695 1526 -2692
rect 1458 -2699 1495 -2695
rect 1458 -2705 1462 -2699
rect 1491 -2705 1495 -2699
rect 2241 -2650 2268 -2647
rect 2241 -2654 2244 -2650
rect 2248 -2654 2261 -2650
rect 2265 -2654 2268 -2650
rect 2241 -2656 2268 -2654
rect 2249 -2661 2253 -2656
rect 2176 -2711 2185 -2710
rect 2069 -2715 2185 -2711
rect 2208 -2711 2212 -2704
rect 2257 -2711 2261 -2701
rect 1514 -2721 1518 -2715
rect 2069 -2716 2178 -2715
rect 2208 -2716 2249 -2711
rect 2257 -2716 2290 -2711
rect 1506 -2722 1533 -2721
rect 1450 -2731 1454 -2725
rect 1483 -2731 1487 -2725
rect 1506 -2726 1507 -2722
rect 1511 -2726 1528 -2722
rect 1532 -2726 1533 -2722
rect 1506 -2727 1533 -2726
rect 1442 -2732 1469 -2731
rect 1442 -2736 1443 -2732
rect 1447 -2736 1464 -2732
rect 1468 -2736 1469 -2732
rect 1442 -2737 1469 -2736
rect 1475 -2732 1502 -2731
rect 1475 -2736 1476 -2732
rect 1480 -2736 1497 -2732
rect 1501 -2736 1502 -2732
rect 1475 -2737 1502 -2736
rect 1464 -2878 1491 -2875
rect 1464 -2882 1467 -2878
rect 1471 -2882 1484 -2878
rect 1488 -2882 1491 -2878
rect 1464 -2884 1491 -2882
rect 1472 -2889 1476 -2884
rect 1358 -2977 1472 -2972
rect 1480 -2981 1484 -2969
rect 1472 -2985 1484 -2981
rect 1472 -2989 1476 -2985
rect 1513 -3015 1540 -3012
rect 1513 -3019 1516 -3015
rect 1520 -3019 1533 -3015
rect 1537 -3019 1540 -3015
rect 1513 -3021 1540 -3019
rect 1521 -3026 1525 -3021
rect 1756 -3034 1783 -3031
rect 1756 -3038 1759 -3034
rect 1763 -3038 1776 -3034
rect 1780 -3038 1783 -3034
rect 1756 -3040 1783 -3038
rect 1341 -3080 1457 -3075
rect 1480 -3076 1484 -3069
rect 1529 -3076 1533 -3066
rect 1764 -3045 1768 -3040
rect 1480 -3081 1521 -3076
rect 1529 -3081 1734 -3076
rect 1480 -3084 1484 -3081
rect 1529 -3084 1533 -3081
rect 1465 -3088 1502 -3084
rect 1465 -3094 1469 -3088
rect 1498 -3094 1502 -3088
rect 1521 -3110 1525 -3104
rect 1513 -3111 1540 -3110
rect 1457 -3120 1461 -3114
rect 1490 -3120 1494 -3114
rect 1513 -3115 1514 -3111
rect 1518 -3115 1535 -3111
rect 1539 -3115 1540 -3111
rect 1513 -3116 1540 -3115
rect 1449 -3121 1476 -3120
rect 1449 -3125 1450 -3121
rect 1454 -3125 1471 -3121
rect 1475 -3125 1476 -3121
rect 1449 -3126 1476 -3125
rect 1482 -3121 1509 -3120
rect 1482 -3125 1483 -3121
rect 1487 -3125 1504 -3121
rect 1508 -3125 1509 -3121
rect 1482 -3126 1509 -3125
rect 1729 -3129 1734 -3081
rect 1747 -3129 1764 -3128
rect 1729 -3133 1764 -3129
rect 1729 -3134 1753 -3133
rect 1772 -3137 1776 -3125
rect 1764 -3141 1776 -3137
rect 1764 -3145 1768 -3141
rect 1805 -3171 1832 -3168
rect 1805 -3175 1808 -3171
rect 1812 -3175 1825 -3171
rect 1829 -3175 1832 -3171
rect 1805 -3177 1832 -3175
rect 1813 -3182 1817 -3177
rect 1458 -3233 1512 -3230
rect 1458 -3237 1461 -3233
rect 1465 -3237 1478 -3233
rect 1482 -3237 1488 -3233
rect 1492 -3237 1505 -3233
rect 1509 -3237 1512 -3233
rect 1458 -3239 1512 -3237
rect 1715 -3236 1749 -3231
rect 1772 -3232 1776 -3225
rect 1821 -3232 1825 -3222
rect 2069 -3232 2074 -2716
rect 2208 -2719 2212 -2716
rect 2257 -2719 2261 -2716
rect 2193 -2723 2230 -2719
rect 2193 -2729 2197 -2723
rect 2226 -2729 2230 -2723
rect 2249 -2745 2253 -2739
rect 2241 -2746 2268 -2745
rect 2185 -2755 2189 -2749
rect 2218 -2755 2222 -2749
rect 2241 -2750 2242 -2746
rect 2246 -2750 2263 -2746
rect 2267 -2750 2268 -2746
rect 2241 -2751 2268 -2750
rect 2177 -2756 2204 -2755
rect 2177 -2760 2178 -2756
rect 2182 -2760 2199 -2756
rect 2203 -2760 2204 -2756
rect 2177 -2761 2204 -2760
rect 2210 -2756 2237 -2755
rect 2210 -2760 2211 -2756
rect 2215 -2760 2232 -2756
rect 2236 -2760 2237 -2756
rect 2210 -2761 2237 -2760
rect 1466 -3244 1470 -3239
rect 1493 -3244 1497 -3239
rect 1474 -3304 1478 -3284
rect 1501 -3304 1505 -3284
rect 1520 -3303 1547 -3300
rect 804 -3434 818 -3430
rect 812 -3435 818 -3434
rect 829 -3435 847 -3430
rect 855 -3435 916 -3430
rect 921 -3309 1463 -3305
rect 1474 -3308 1515 -3304
rect 921 -3310 1466 -3309
rect 325 -3446 326 -3441
rect 331 -3446 804 -3441
rect 812 -3449 816 -3435
rect 855 -3438 859 -3435
rect 847 -3464 851 -3458
rect 839 -3465 866 -3464
rect 839 -3469 840 -3465
rect 844 -3469 861 -3465
rect 865 -3469 866 -3465
rect 839 -3470 866 -3469
rect 804 -3495 808 -3489
rect 796 -3496 823 -3495
rect 796 -3500 797 -3496
rect 801 -3500 818 -3496
rect 822 -3500 823 -3496
rect 796 -3501 823 -3500
rect 794 -3566 848 -3563
rect 794 -3570 797 -3566
rect 801 -3570 814 -3566
rect 818 -3570 824 -3566
rect 828 -3570 841 -3566
rect 845 -3570 848 -3566
rect 794 -3572 848 -3570
rect 802 -3577 806 -3572
rect 829 -3577 833 -3572
rect 810 -3637 814 -3617
rect 837 -3637 841 -3617
rect 856 -3636 883 -3633
rect 810 -3641 851 -3637
rect 298 -3647 299 -3642
rect 304 -3647 802 -3642
rect 829 -3651 833 -3641
rect 821 -3697 825 -3691
rect 846 -3697 851 -3641
rect 856 -3640 859 -3636
rect 863 -3640 876 -3636
rect 880 -3640 883 -3636
rect 856 -3642 883 -3640
rect 864 -3647 868 -3642
rect 872 -3697 876 -3687
rect 921 -3697 926 -3310
rect 1458 -3314 1466 -3310
rect 1458 -3315 1463 -3314
rect 1493 -3318 1497 -3308
rect 1118 -3365 1172 -3362
rect 1118 -3369 1121 -3365
rect 1125 -3369 1138 -3365
rect 1142 -3369 1148 -3365
rect 1152 -3369 1165 -3365
rect 1169 -3369 1172 -3365
rect 1485 -3364 1489 -3358
rect 1510 -3364 1515 -3308
rect 1520 -3307 1523 -3303
rect 1527 -3307 1540 -3303
rect 1544 -3307 1547 -3303
rect 1520 -3309 1547 -3307
rect 1528 -3314 1532 -3309
rect 1536 -3364 1540 -3354
rect 1715 -3364 1720 -3236
rect 1772 -3237 1813 -3232
rect 1821 -3237 2074 -3232
rect 1772 -3240 1776 -3237
rect 1821 -3240 1825 -3237
rect 1757 -3244 1794 -3240
rect 1757 -3250 1761 -3244
rect 1790 -3250 1794 -3244
rect 1813 -3266 1817 -3260
rect 1805 -3267 1832 -3266
rect 1749 -3276 1753 -3270
rect 1782 -3276 1786 -3270
rect 1805 -3271 1806 -3267
rect 1810 -3271 1827 -3267
rect 1831 -3271 1832 -3267
rect 1805 -3272 1832 -3271
rect 1741 -3277 1768 -3276
rect 1741 -3281 1742 -3277
rect 1746 -3281 1763 -3277
rect 1767 -3281 1768 -3277
rect 1741 -3282 1768 -3281
rect 1774 -3277 1801 -3276
rect 1774 -3281 1775 -3277
rect 1779 -3281 1796 -3277
rect 1800 -3281 1801 -3277
rect 1774 -3282 1801 -3281
rect 1485 -3368 1499 -3364
rect 1118 -3371 1172 -3369
rect 1493 -3369 1499 -3368
rect 1510 -3369 1528 -3364
rect 1536 -3369 1720 -3364
rect 1126 -3376 1130 -3371
rect 1153 -3376 1157 -3371
rect 1134 -3436 1138 -3416
rect 1161 -3436 1165 -3416
rect 1261 -3380 1485 -3375
rect 1180 -3435 1207 -3432
rect 1119 -3441 1124 -3439
rect 1134 -3440 1175 -3436
rect 1119 -3443 1126 -3441
rect 821 -3701 835 -3697
rect 829 -3702 835 -3701
rect 846 -3702 864 -3697
rect 872 -3702 926 -3697
rect 1006 -3446 1126 -3443
rect 1006 -3448 1124 -3446
rect 307 -3713 308 -3708
rect 313 -3713 821 -3708
rect 829 -3716 833 -3702
rect 872 -3705 876 -3702
rect 864 -3731 868 -3725
rect 856 -3732 883 -3731
rect 856 -3736 857 -3732
rect 861 -3736 878 -3732
rect 882 -3736 883 -3732
rect 856 -3737 883 -3736
rect 821 -3762 825 -3756
rect 813 -3763 840 -3762
rect 813 -3767 814 -3763
rect 818 -3767 835 -3763
rect 839 -3767 840 -3763
rect 813 -3768 840 -3767
rect 782 -3815 836 -3812
rect 782 -3819 785 -3815
rect 789 -3819 802 -3815
rect 806 -3819 812 -3815
rect 816 -3819 829 -3815
rect 833 -3819 836 -3815
rect 782 -3821 836 -3819
rect 790 -3826 794 -3821
rect 817 -3826 821 -3821
rect 798 -3886 802 -3866
rect 825 -3886 829 -3866
rect 844 -3885 871 -3882
rect 798 -3890 839 -3886
rect 325 -3896 326 -3891
rect 331 -3896 790 -3891
rect 817 -3900 821 -3890
rect 809 -3946 813 -3940
rect 834 -3946 839 -3890
rect 844 -3889 847 -3885
rect 851 -3889 864 -3885
rect 868 -3889 871 -3885
rect 844 -3891 871 -3889
rect 852 -3896 856 -3891
rect 860 -3946 864 -3936
rect 1006 -3946 1011 -3448
rect 1119 -3450 1124 -3448
rect 1153 -3450 1157 -3440
rect 1145 -3496 1149 -3490
rect 1170 -3496 1175 -3440
rect 1180 -3439 1183 -3435
rect 1187 -3439 1200 -3435
rect 1204 -3439 1207 -3435
rect 1180 -3441 1207 -3439
rect 1188 -3446 1192 -3441
rect 1196 -3496 1200 -3486
rect 1261 -3495 1266 -3380
rect 1493 -3383 1497 -3369
rect 1536 -3372 1540 -3369
rect 1528 -3398 1532 -3392
rect 1520 -3399 1547 -3398
rect 1520 -3403 1521 -3399
rect 1525 -3403 1542 -3399
rect 1546 -3403 1547 -3399
rect 1520 -3404 1547 -3403
rect 1485 -3429 1489 -3423
rect 1477 -3430 1504 -3429
rect 1477 -3434 1478 -3430
rect 1482 -3434 1499 -3430
rect 1503 -3434 1504 -3430
rect 1477 -3435 1504 -3434
rect 1206 -3496 1266 -3495
rect 1145 -3500 1159 -3496
rect 1153 -3501 1159 -3500
rect 1170 -3501 1188 -3496
rect 1196 -3500 1266 -3496
rect 1196 -3501 1209 -3500
rect 809 -3950 823 -3946
rect 817 -3951 823 -3950
rect 834 -3951 852 -3946
rect 860 -3951 1011 -3946
rect 1052 -3512 1145 -3507
rect 343 -3962 344 -3957
rect 349 -3962 809 -3957
rect 817 -3965 821 -3951
rect 860 -3954 864 -3951
rect 852 -3980 856 -3974
rect 844 -3981 871 -3980
rect 844 -3985 845 -3981
rect 849 -3985 866 -3981
rect 870 -3985 871 -3981
rect 844 -3986 871 -3985
rect 809 -4011 813 -4005
rect 801 -4012 828 -4011
rect 801 -4016 802 -4012
rect 806 -4016 823 -4012
rect 827 -4016 828 -4012
rect 801 -4017 828 -4016
rect 1052 -4026 1057 -3512
rect 1153 -3515 1157 -3501
rect 1196 -3504 1200 -3501
rect 1188 -3530 1192 -3524
rect 1180 -3531 1207 -3530
rect 1180 -3535 1181 -3531
rect 1185 -3535 1202 -3531
rect 1206 -3535 1207 -3531
rect 1180 -3536 1207 -3535
rect 1145 -3561 1149 -3555
rect 1137 -3562 1164 -3561
rect 1137 -3566 1138 -3562
rect 1142 -3566 1159 -3562
rect 1163 -3566 1164 -3562
rect 1137 -3567 1164 -3566
rect 361 -4031 362 -4026
rect 367 -4031 1057 -4026
<< m2contact >>
rect 299 26 304 31
rect 308 -22 313 -17
rect 14 -176 19 -171
rect 308 -218 313 -213
rect 299 -284 304 -279
rect 101 -377 107 -372
rect 317 -432 322 -427
rect 326 -461 331 -456
rect 335 -864 340 -859
rect 317 -888 322 -883
rect 2 -962 7 -957
rect 326 -1004 331 -999
rect 299 -1133 304 -1128
rect 308 -1145 313 -1140
rect 89 -1163 95 -1158
rect 335 -1218 340 -1213
rect 326 -1271 331 -1266
rect 344 -1305 349 -1299
rect 353 -1319 358 -1314
rect 344 -1425 349 -1420
rect 335 -1491 340 -1486
rect 11 -1622 16 -1617
rect 344 -1664 349 -1659
rect 344 -1708 349 -1703
rect 326 -1774 331 -1769
rect 98 -1823 104 -1818
rect 317 -1845 322 -1840
rect 353 -1878 358 -1873
rect 299 -1979 304 -1974
rect 308 -2045 313 -2040
rect 344 -2228 349 -2223
rect 326 -2294 331 -2289
rect 362 -2383 367 -2378
rect 8 -2497 13 -2492
rect 362 -2539 367 -2534
rect 95 -2698 101 -2693
rect 353 -2770 358 -2765
rect 362 -2779 367 -2774
rect 362 -2860 367 -2855
rect 344 -2926 349 -2921
rect 335 -3000 340 -2995
rect 362 -3131 367 -3126
rect 344 -3197 349 -3192
rect 317 -3380 322 -3375
rect 326 -3446 331 -3441
rect 299 -3647 304 -3642
rect 308 -3713 313 -3708
rect 326 -3896 331 -3891
rect 344 -3962 349 -3957
rect 362 -4031 367 -4026
<< metal2 >>
rect 14 -372 19 -176
rect 299 -279 304 26
rect 14 -377 101 -372
rect 2 -1158 7 -962
rect 299 -1128 304 -284
rect 2 -1163 89 -1158
rect 11 -1818 16 -1622
rect 11 -1823 98 -1818
rect 299 -1974 304 -1133
rect 8 -2693 13 -2497
rect 8 -2698 95 -2693
rect 299 -3642 304 -1979
rect 299 -4035 304 -3647
rect 308 -213 313 -22
rect 308 -1140 313 -218
rect 308 -2040 313 -1145
rect 308 -3708 313 -2045
rect 308 -4036 313 -3713
rect 317 -883 322 -432
rect 317 -1840 322 -888
rect 317 -3375 322 -1845
rect 317 -4032 322 -3380
rect 326 -999 331 -461
rect 326 -1266 331 -1004
rect 326 -1769 331 -1271
rect 326 -2289 331 -1774
rect 326 -3441 331 -2294
rect 326 -3891 331 -3446
rect 326 -4034 331 -3896
rect 335 -1213 340 -864
rect 335 -1486 340 -1218
rect 335 -2995 340 -1491
rect 335 -4033 340 -3000
rect 344 -1420 349 -1305
rect 344 -1659 349 -1425
rect 344 -1703 349 -1664
rect 344 -2223 349 -1708
rect 344 -2921 349 -2228
rect 344 -3192 349 -2926
rect 344 -3957 349 -3197
rect 344 -4033 349 -3962
rect 353 -1873 358 -1319
rect 353 -2765 358 -1878
rect 353 -4034 358 -2770
rect 362 -2378 367 -2373
rect 362 -2534 367 -2383
rect 362 -2774 367 -2539
rect 362 -2855 367 -2779
rect 362 -3126 367 -2860
rect 362 -4026 367 -3131
rect 362 -4034 367 -4031
<< labels >>
rlabel metal1 207 -243 207 -243 7 vdd
rlabel metal1 111 -243 111 -243 3 gnd
rlabel metal1 207 -192 207 -192 7 vdd
rlabel metal1 111 -192 111 -192 3 gnd
rlabel metal1 259 -250 259 -250 1 gnd
rlabel metal1 259 -154 259 -154 5 vdd
rlabel metal1 176 -298 176 -298 5 vdd
rlabel metal1 203 -298 203 -298 5 vdd
rlabel metal1 195 -495 195 -495 1 gnd
rlabel metal1 238 -368 238 -368 5 vdd
rlabel metal1 238 -464 238 -464 1 gnd
rlabel metal1 -10 -174 -10 -174 1 A0
rlabel metal1 -13 -221 -13 -221 1 B0
rlabel metal1 292 -430 292 -430 1 G0
rlabel metal1 2095 -1072 2095 -1072 7 vdd
rlabel metal1 1999 -1072 1999 -1072 3 gnd
rlabel metal1 2095 -1021 2095 -1021 7 vdd
rlabel metal1 1999 -1021 1999 -1021 3 gnd
rlabel metal1 2147 -1079 2147 -1079 1 gnd
rlabel metal1 2147 -983 2147 -983 5 vdd
rlabel metal1 2093 -1780 2093 -1780 7 vdd
rlabel metal1 1997 -1780 1997 -1780 3 gnd
rlabel metal1 2093 -1729 2093 -1729 7 vdd
rlabel metal1 1997 -1729 1997 -1729 3 gnd
rlabel metal1 2145 -1787 2145 -1787 1 gnd
rlabel metal1 2145 -1691 2145 -1691 5 vdd
rlabel metal1 1776 -1859 1776 -1859 1 gnd
rlabel metal1 1776 -1763 1776 -1763 5 vdd
rlabel metal1 1745 -1869 1745 -1869 1 gnd
rlabel metal1 1712 -1869 1712 -1869 1 gnd
rlabel metal1 1727 -1626 1727 -1626 5 vdd
rlabel metal1 1479 -1706 1479 -1706 1 gnd
rlabel metal1 1479 -1610 1479 -1610 5 vdd
rlabel metal1 1448 -1716 1448 -1716 1 gnd
rlabel metal1 1415 -1716 1415 -1716 1 gnd
rlabel metal1 1430 -1473 1430 -1473 5 vdd
rlabel metal1 1490 -2006 1490 -2006 1 gnd
rlabel metal1 1490 -1910 1490 -1910 5 vdd
rlabel metal1 1459 -2016 1459 -2016 1 gnd
rlabel metal1 1426 -2016 1426 -2016 1 gnd
rlabel metal1 1441 -1773 1441 -1773 5 vdd
rlabel metal1 1078 -1646 1078 -1646 5 vdd
rlabel metal1 1035 -1773 1035 -1773 1 gnd
rlabel metal1 1043 -1576 1043 -1576 5 vdd
rlabel metal1 1016 -1576 1016 -1576 5 vdd
rlabel metal1 1087 -1953 1087 -1953 1 gnd
rlabel metal1 1087 -1857 1087 -1857 5 vdd
rlabel metal1 1044 -1984 1044 -1984 1 gnd
rlabel metal1 1052 -1787 1052 -1787 5 vdd
rlabel metal1 1025 -1787 1025 -1787 5 vdd
rlabel metal1 1683 -42 1683 -42 7 vdd
rlabel metal1 1587 -42 1587 -42 3 gnd
rlabel metal1 1683 9 1683 9 7 vdd
rlabel metal1 1587 9 1587 9 3 gnd
rlabel metal1 1735 -49 1735 -49 1 gnd
rlabel metal1 1735 47 1735 47 5 vdd
rlabel metal1 1678 -262 1678 -262 7 vdd
rlabel metal1 1582 -262 1582 -262 3 gnd
rlabel metal1 1678 -211 1678 -211 7 vdd
rlabel metal1 1582 -211 1582 -211 3 gnd
rlabel metal1 1730 -269 1730 -269 1 gnd
rlabel metal1 1730 -173 1730 -173 5 vdd
rlabel metal1 1104 -54 1104 -54 5 vdd
rlabel metal1 1089 -297 1089 -297 1 gnd
rlabel metal1 1122 -297 1122 -297 1 gnd
rlabel metal1 1153 -191 1153 -191 5 vdd
rlabel metal1 1153 -287 1153 -287 1 gnd
rlabel metal1 1793 -1011 1793 -1011 1 gnd
rlabel metal1 1793 -915 1793 -915 5 vdd
rlabel metal1 1762 -1021 1762 -1021 1 gnd
rlabel metal1 1729 -1021 1729 -1021 1 gnd
rlabel metal1 1744 -778 1744 -778 5 vdd
rlabel metal1 1542 -1009 1542 -1009 1 gnd
rlabel metal1 1542 -913 1542 -913 5 vdd
rlabel metal1 1511 -1019 1511 -1019 1 gnd
rlabel metal1 1478 -1019 1478 -1019 1 gnd
rlabel metal1 1493 -776 1493 -776 5 vdd
rlabel metal1 1156 -975 1156 -975 1 gnd
rlabel metal1 1156 -879 1156 -879 5 vdd
rlabel metal1 1113 -1006 1113 -1006 1 gnd
rlabel metal1 1121 -809 1121 -809 5 vdd
rlabel metal1 1094 -809 1094 -809 5 vdd
rlabel metal1 1079 -1220 1079 -1220 1 gnd
rlabel metal1 1079 -1124 1079 -1124 5 vdd
rlabel metal1 1036 -1251 1036 -1251 1 gnd
rlabel metal1 1044 -1054 1044 -1054 5 vdd
rlabel metal1 1017 -1054 1017 -1054 5 vdd
rlabel metal1 1297 -1220 1297 -1220 1 gnd
rlabel metal1 1297 -1124 1297 -1124 5 vdd
rlabel metal1 1254 -1251 1254 -1251 1 gnd
rlabel metal1 1262 -1054 1262 -1054 5 vdd
rlabel metal1 1235 -1054 1235 -1054 5 vdd
rlabel metal1 838 -2066 838 -2066 1 gnd
rlabel metal1 838 -1970 838 -1970 5 vdd
rlabel metal1 795 -2097 795 -2097 1 gnd
rlabel metal1 803 -1900 803 -1900 5 vdd
rlabel metal1 776 -1900 776 -1900 5 vdd
rlabel metal1 842 -1795 842 -1795 1 gnd
rlabel metal1 842 -1699 842 -1699 5 vdd
rlabel metal1 799 -1826 799 -1826 1 gnd
rlabel metal1 807 -1629 807 -1629 5 vdd
rlabel metal1 780 -1629 780 -1629 5 vdd
rlabel metal1 841 -1512 841 -1512 1 gnd
rlabel metal1 841 -1416 841 -1416 5 vdd
rlabel metal1 798 -1543 798 -1543 1 gnd
rlabel metal1 806 -1346 806 -1346 5 vdd
rlabel metal1 779 -1346 779 -1346 5 vdd
rlabel metal1 826 -2315 826 -2315 1 gnd
rlabel metal1 826 -2219 826 -2219 5 vdd
rlabel metal1 791 -2149 791 -2149 5 vdd
rlabel metal1 764 -2149 764 -2149 5 vdd
rlabel metal1 783 -2346 783 -2346 1 gnd
rlabel metal1 1519 -2724 1519 -2724 1 gnd
rlabel metal1 1519 -2628 1519 -2628 5 vdd
rlabel metal1 1488 -2734 1488 -2734 1 gnd
rlabel metal1 1455 -2734 1455 -2734 1 gnd
rlabel metal1 1470 -2491 1470 -2491 5 vdd
rlabel metal1 1526 -3113 1526 -3113 1 gnd
rlabel metal1 1526 -3017 1526 -3017 5 vdd
rlabel metal1 1495 -3123 1495 -3123 1 gnd
rlabel metal1 1462 -3123 1462 -3123 1 gnd
rlabel metal1 1477 -2880 1477 -2880 5 vdd
rlabel metal1 1818 -3269 1818 -3269 1 gnd
rlabel metal1 1818 -3173 1818 -3173 5 vdd
rlabel metal1 1787 -3279 1787 -3279 1 gnd
rlabel metal1 1754 -3279 1754 -3279 1 gnd
rlabel metal1 1769 -3036 1769 -3036 5 vdd
rlabel metal1 2254 -2748 2254 -2748 1 gnd
rlabel metal1 2254 -2652 2254 -2652 5 vdd
rlabel metal1 2223 -2758 2223 -2758 1 gnd
rlabel metal1 2190 -2758 2190 -2758 1 gnd
rlabel metal1 2205 -2515 2205 -2515 5 vdd
rlabel metal1 1078 -1742 1078 -1742 1 gnd
rlabel metal1 864 -3218 864 -3218 1 gnd
rlabel metal1 864 -3122 864 -3122 5 vdd
rlabel metal1 821 -3249 821 -3249 1 gnd
rlabel metal1 829 -3052 829 -3052 5 vdd
rlabel metal1 802 -3052 802 -3052 5 vdd
rlabel metal1 868 -2947 868 -2947 1 gnd
rlabel metal1 868 -2851 868 -2851 5 vdd
rlabel metal1 825 -2978 825 -2978 1 gnd
rlabel metal1 833 -2781 833 -2781 5 vdd
rlabel metal1 806 -2781 806 -2781 5 vdd
rlabel metal1 867 -2664 867 -2664 1 gnd
rlabel metal1 867 -2568 867 -2568 5 vdd
rlabel metal1 824 -2695 824 -2695 1 gnd
rlabel metal1 832 -2498 832 -2498 5 vdd
rlabel metal1 805 -2498 805 -2498 5 vdd
rlabel metal1 852 -3467 852 -3467 1 gnd
rlabel metal1 852 -3371 852 -3371 5 vdd
rlabel metal1 817 -3301 817 -3301 5 vdd
rlabel metal1 790 -3301 790 -3301 5 vdd
rlabel metal1 809 -3498 809 -3498 1 gnd
rlabel metal1 1203 -2999 1203 -2999 1 gnd
rlabel metal1 1203 -2903 1203 -2903 5 vdd
rlabel metal1 1160 -3030 1160 -3030 1 gnd
rlabel metal1 1168 -2833 1168 -2833 5 vdd
rlabel metal1 1141 -2833 1141 -2833 5 vdd
rlabel metal1 1202 -2716 1202 -2716 1 gnd
rlabel metal1 1202 -2620 1202 -2620 5 vdd
rlabel metal1 1159 -2747 1159 -2747 1 gnd
rlabel metal1 1167 -2550 1167 -2550 5 vdd
rlabel metal1 1140 -2550 1140 -2550 5 vdd
rlabel metal1 869 -3734 869 -3734 1 gnd
rlabel metal1 869 -3638 869 -3638 5 vdd
rlabel metal1 826 -3765 826 -3765 1 gnd
rlabel metal1 834 -3568 834 -3568 5 vdd
rlabel metal1 807 -3568 807 -3568 5 vdd
rlabel metal1 857 -3983 857 -3983 1 gnd
rlabel metal1 857 -3887 857 -3887 5 vdd
rlabel metal1 822 -3817 822 -3817 5 vdd
rlabel metal1 795 -3817 795 -3817 5 vdd
rlabel metal1 814 -4014 814 -4014 1 gnd
rlabel metal1 287 -216 287 -216 1 P0
rlabel metal1 796 -305 796 -305 1 gnd
rlabel metal1 796 -209 796 -209 5 vdd
rlabel metal1 753 -336 753 -336 1 gnd
rlabel metal1 761 -139 761 -139 5 vdd
rlabel metal1 734 -139 734 -139 5 vdd
rlabel metal1 204 -1689 204 -1689 7 vdd
rlabel metal1 108 -1689 108 -1689 3 gnd
rlabel metal1 204 -1638 204 -1638 7 vdd
rlabel metal1 108 -1638 108 -1638 3 gnd
rlabel metal1 256 -1696 256 -1696 1 gnd
rlabel metal1 256 -1600 256 -1600 5 vdd
rlabel metal1 173 -1744 173 -1744 5 vdd
rlabel metal1 200 -1744 200 -1744 5 vdd
rlabel metal1 192 -1941 192 -1941 1 gnd
rlabel metal1 235 -1814 235 -1814 5 vdd
rlabel metal1 235 -1910 235 -1910 1 gnd
rlabel metal1 -15 -1620 -15 -1620 1 A2
rlabel metal1 -17 -1667 -17 -1667 1 B2
rlabel metal1 290 -1662 290 -1662 1 P2
rlabel metal1 287 -1876 287 -1876 1 G2
rlabel metal1 195 -1029 195 -1029 7 vdd
rlabel metal1 99 -1029 99 -1029 3 gnd
rlabel metal1 195 -978 195 -978 7 vdd
rlabel metal1 99 -978 99 -978 3 gnd
rlabel metal1 247 -1036 247 -1036 1 gnd
rlabel metal1 247 -940 247 -940 5 vdd
rlabel metal1 164 -1084 164 -1084 5 vdd
rlabel metal1 191 -1084 191 -1084 5 vdd
rlabel metal1 183 -1281 183 -1281 1 gnd
rlabel metal1 226 -1154 226 -1154 5 vdd
rlabel metal1 226 -1250 226 -1250 1 gnd
rlabel metal1 -27 -960 -27 -960 1 A1
rlabel metal1 -23 -1007 -23 -1007 1 B1
rlabel metal1 281 -1002 281 -1002 1 P1
rlabel metal1 281 -1216 281 -1216 1 G1
rlabel metal1 201 -2564 201 -2564 7 vdd
rlabel metal1 105 -2564 105 -2564 3 gnd
rlabel metal1 201 -2513 201 -2513 7 vdd
rlabel metal1 105 -2513 105 -2513 3 gnd
rlabel metal1 253 -2571 253 -2571 1 gnd
rlabel metal1 253 -2475 253 -2475 5 vdd
rlabel metal1 170 -2619 170 -2619 5 vdd
rlabel metal1 197 -2619 197 -2619 5 vdd
rlabel metal1 189 -2816 189 -2816 1 gnd
rlabel metal1 232 -2689 232 -2689 5 vdd
rlabel metal1 232 -2785 232 -2785 1 gnd
rlabel metal1 -21 -2494 -21 -2494 1 A3
rlabel metal1 -18 -2542 -18 -2542 1 B3
rlabel metal1 287 -2537 287 -2537 1 P3
rlabel metal1 284 -2751 284 -2751 1 G3
rlabel metal1 1173 -251 1173 -251 1 c1
rlabel metal1 -14 28 -14 28 1 c0
rlabel metal1 1533 -3401 1533 -3401 1 gnd
rlabel metal1 1533 -3305 1533 -3305 5 vdd
rlabel metal1 1490 -3432 1490 -3432 1 gnd
rlabel metal1 1498 -3235 1498 -3235 5 vdd
rlabel metal1 1471 -3235 1471 -3235 5 vdd
rlabel metal1 1193 -3533 1193 -3533 1 gnd
rlabel metal1 1193 -3437 1193 -3437 5 vdd
rlabel metal1 1158 -3367 1158 -3367 5 vdd
rlabel metal1 1131 -3367 1131 -3367 5 vdd
rlabel metal1 1150 -3564 1150 -3564 1 gnd
rlabel metal1 -3492 -1263 -3492 -1263 7 vdd
rlabel metal1 -3588 -1263 -3588 -1263 3 gnd
rlabel metal1 -3492 -1212 -3492 -1212 7 vdd
rlabel metal1 -3588 -1212 -3588 -1212 3 gnd
rlabel metal1 -3440 -1270 -3440 -1270 1 gnd
rlabel metal1 -3440 -1174 -3440 -1174 5 vdd
rlabel metal1 -3113 -1325 -3113 -1325 1 gnd
rlabel metal1 -3113 -1229 -3113 -1229 5 vdd
rlabel metal1 -3156 -1356 -3156 -1356 1 gnd
rlabel metal1 -3148 -1159 -3148 -1159 5 vdd
rlabel metal1 -3175 -1159 -3175 -1159 5 vdd
rlabel metal1 -3235 -1380 -3235 -1380 1 gnd
rlabel metal1 -3235 -1284 -3235 -1284 5 vdd
rlabel metal1 -3266 -1390 -3266 -1390 1 gnd
rlabel metal1 -3299 -1390 -3299 -1390 1 gnd
rlabel metal1 -3284 -1147 -3284 -1147 5 vdd
rlabel metal1 -3349 -1286 -3349 -1286 1 gnd
rlabel metal1 -3349 -1190 -3349 -1190 5 vdd
rlabel metal1 1769 -15 1769 -15 1 S0
rlabel metal1 1759 -234 1759 -234 1 S1
rlabel metal1 2159 -1045 2159 -1045 1 S2
rlabel metal1 2156 -1753 2156 -1753 1 S3
rlabel metal1 2266 -2713 2266 -2713 7 S4
rlabel metal1 2266 -2713 2266 -2713 7 Cout
rlabel metal1 2286 -2714 2286 -2713 7 Cout
<< end >>
