magic
tech scmos
timestamp 1731695926
<< nwell >>
rect -118 291 -56 318
rect -22 286 5 348
rect 69 270 96 332
rect -118 240 -56 267
rect 134 173 161 375
rect 243 301 297 363
rect 183 176 210 238
rect 305 231 332 293
<< ntransistor >>
rect -148 303 -128 305
rect -45 291 -43 311
rect -45 258 -43 278
rect -9 256 -7 276
rect -148 252 -128 254
rect 82 240 84 260
rect 275 235 277 275
rect 275 170 277 210
rect 318 201 320 221
rect 132 136 134 156
rect 165 136 167 156
rect 196 146 198 166
<< ptransistor >>
rect -110 303 -70 305
rect -9 294 -7 334
rect 82 278 84 318
rect 147 281 149 361
rect 256 309 258 349
rect 283 309 285 349
rect -110 252 -70 254
rect 147 181 149 261
rect 196 184 198 224
rect 318 239 320 279
<< ndiffusion >>
rect -148 305 -128 306
rect -148 302 -128 303
rect -46 291 -45 311
rect -43 291 -42 311
rect -148 254 -128 255
rect -46 258 -45 278
rect -43 258 -42 278
rect -10 256 -9 276
rect -7 256 -6 276
rect -148 251 -128 252
rect 81 240 82 260
rect 84 240 85 260
rect 274 235 275 275
rect 277 235 278 275
rect 274 170 275 210
rect 277 170 278 210
rect 317 201 318 221
rect 320 201 321 221
rect 131 136 132 156
rect 134 136 135 156
rect 164 136 165 156
rect 167 136 168 156
rect 195 146 196 166
rect 198 146 199 166
<< pdiffusion >>
rect -110 305 -70 306
rect -110 302 -70 303
rect -10 294 -9 334
rect -7 294 -6 334
rect 81 278 82 318
rect 84 278 85 318
rect 146 281 147 361
rect 149 281 150 361
rect 255 309 256 349
rect 258 309 259 349
rect 282 309 283 349
rect 285 309 286 349
rect -110 254 -70 255
rect -110 251 -70 252
rect 146 181 147 261
rect 149 181 150 261
rect 195 184 196 224
rect 198 184 199 224
rect 317 239 318 279
rect 320 239 321 279
<< ndcontact >>
rect -148 306 -128 310
rect -148 298 -128 302
rect -50 291 -46 311
rect -42 291 -38 311
rect -148 255 -128 259
rect -50 258 -46 278
rect -42 258 -38 278
rect -14 256 -10 276
rect -6 256 -2 276
rect -148 247 -128 251
rect 77 240 81 260
rect 85 240 89 260
rect 270 235 274 275
rect 278 235 282 275
rect 270 170 274 210
rect 278 170 282 210
rect 313 201 317 221
rect 321 201 325 221
rect 127 136 131 156
rect 135 136 139 156
rect 160 136 164 156
rect 168 136 172 156
rect 191 146 195 166
rect 199 146 203 166
<< pdcontact >>
rect -110 306 -70 310
rect -110 298 -70 302
rect -14 294 -10 334
rect -6 294 -2 334
rect -110 255 -70 259
rect 77 278 81 318
rect 85 278 89 318
rect 142 281 146 361
rect 150 281 154 361
rect 251 309 255 349
rect 259 309 263 349
rect 278 309 282 349
rect 286 309 290 349
rect -110 247 -70 251
rect 142 181 146 261
rect 150 181 154 261
rect 191 184 195 224
rect 199 184 203 224
rect 313 239 317 279
rect 321 239 325 279
<< psubstratepcontact >>
rect -159 313 -155 317
rect -159 292 -155 296
rect -159 262 -155 266
rect -159 241 -155 245
rect -21 245 -17 249
rect 0 245 4 249
rect 70 229 74 233
rect 91 229 95 233
rect 306 190 310 194
rect 327 190 331 194
rect 263 159 267 163
rect 284 159 288 163
rect 184 135 188 139
rect 205 135 209 139
rect 120 125 124 129
rect 141 125 145 129
rect 153 125 157 129
rect 174 125 178 129
<< nsubstratencontact >>
rect 137 368 141 372
rect 154 368 158 372
rect -19 341 -15 345
rect -2 341 2 345
rect -63 311 -59 315
rect -63 294 -59 298
rect 72 325 76 329
rect 89 325 93 329
rect -63 260 -59 264
rect 246 356 250 360
rect 263 356 267 360
rect 273 356 277 360
rect 290 356 294 360
rect -63 243 -59 247
rect 186 231 190 235
rect 203 231 207 235
rect 308 286 312 290
rect 325 286 329 290
<< polysilicon >>
rect 147 361 149 364
rect -125 333 -43 335
rect -9 334 -7 337
rect -45 311 -43 333
rect -151 303 -148 305
rect -128 303 -110 305
rect -70 303 -67 305
rect 82 318 84 321
rect -45 288 -43 291
rect -125 281 -43 283
rect -45 278 -43 281
rect -9 276 -7 294
rect 256 349 258 352
rect 283 349 285 352
rect -45 255 -43 258
rect 82 260 84 278
rect 147 275 149 281
rect 256 281 258 309
rect 283 297 285 309
rect 283 295 293 297
rect 256 279 277 281
rect 275 275 277 279
rect 147 273 167 275
rect 147 261 149 264
rect -151 252 -148 254
rect -128 252 -110 254
rect -70 252 -67 254
rect -9 253 -7 256
rect 82 237 84 240
rect 147 175 149 181
rect 132 173 149 175
rect 132 156 134 173
rect 165 156 167 273
rect 275 231 277 235
rect 196 224 198 227
rect 291 218 293 295
rect 318 279 320 282
rect 318 221 320 239
rect 275 216 293 218
rect 275 210 277 216
rect 196 166 198 184
rect 318 198 320 201
rect 275 167 277 170
rect 196 143 198 146
rect 132 133 134 136
rect 165 133 167 136
<< polycontact >>
rect -125 328 -120 333
rect -125 305 -120 310
rect -125 283 -120 288
rect -14 279 -9 284
rect -125 254 -120 259
rect 77 263 82 268
rect 142 273 147 278
rect 251 279 256 284
rect 127 170 132 175
rect 313 224 318 229
rect 270 213 275 218
rect 191 169 196 174
<< metal1 >>
rect 134 372 161 375
rect 134 368 137 372
rect 141 368 154 372
rect 158 368 161 372
rect 134 366 161 368
rect 142 361 146 366
rect -22 345 5 348
rect -22 341 -19 345
rect -15 341 -2 345
rect 2 341 5 345
rect -22 339 5 341
rect -14 334 -10 339
rect -125 326 -120 328
rect -160 321 -120 326
rect -160 317 -154 318
rect -160 313 -159 317
rect -155 313 -154 317
rect -160 310 -154 313
rect -125 310 -120 321
rect -65 315 -56 318
rect -65 311 -63 315
rect -59 311 -56 315
rect -42 311 -29 314
rect -65 310 -56 311
rect -160 306 -148 310
rect -160 296 -154 306
rect -70 306 -56 310
rect -128 298 -110 302
rect -65 298 -56 306
rect -160 292 -159 296
rect -155 292 -154 296
rect -160 291 -154 292
rect -125 288 -120 298
rect -65 294 -63 298
rect -59 294 -56 298
rect -65 291 -56 294
rect -50 288 -46 291
rect -96 284 -46 288
rect -96 279 -92 284
rect -160 274 -92 279
rect -42 278 -38 291
rect -35 284 -29 311
rect 69 329 96 332
rect 69 325 72 329
rect 76 325 89 329
rect 93 325 96 329
rect 69 323 96 325
rect -6 284 -2 294
rect 77 318 81 323
rect -35 279 -14 284
rect -6 279 5 284
rect -160 266 -154 267
rect -160 262 -159 266
rect -155 262 -154 266
rect -160 259 -154 262
rect -125 259 -120 274
rect -65 264 -56 267
rect -65 260 -63 264
rect -59 260 -56 264
rect -65 259 -56 260
rect -160 255 -148 259
rect -160 245 -154 255
rect -70 255 -56 259
rect -128 247 -110 251
rect -65 247 -56 255
rect -160 241 -159 245
rect -155 241 -154 245
rect -160 240 -154 241
rect -125 227 -120 247
rect -65 243 -63 247
rect -59 243 -56 247
rect -65 240 -56 243
rect -6 276 -2 279
rect 243 360 297 363
rect 243 356 246 360
rect 250 356 263 360
rect 267 356 273 360
rect 277 356 290 360
rect 294 356 297 360
rect 243 354 297 356
rect 251 349 255 354
rect 278 349 282 354
rect 259 289 263 309
rect 286 289 290 309
rect 305 290 332 293
rect 259 285 300 289
rect -50 227 -46 258
rect 85 268 89 278
rect 125 273 142 278
rect 150 269 154 281
rect 244 279 251 284
rect 278 275 282 285
rect 69 263 77 268
rect 85 263 98 268
rect 142 265 154 269
rect 85 260 89 263
rect -14 250 -10 256
rect -22 249 5 250
rect -22 245 -21 249
rect -17 245 0 249
rect 4 245 5 249
rect -22 244 5 245
rect 142 261 146 265
rect 77 234 81 240
rect 69 233 96 234
rect 69 229 70 233
rect 74 229 91 233
rect 95 229 96 233
rect 69 228 96 229
rect -125 224 -46 227
rect 183 235 210 238
rect 183 231 186 235
rect 190 231 203 235
rect 207 231 210 235
rect 183 229 210 231
rect 270 229 274 235
rect 295 229 300 285
rect 305 286 308 290
rect 312 286 325 290
rect 329 286 332 290
rect 305 284 332 286
rect 313 279 317 284
rect 321 229 325 239
rect 191 224 195 229
rect 270 225 284 229
rect 278 224 284 225
rect 295 224 313 229
rect 321 224 334 229
rect 244 213 270 218
rect 278 210 282 224
rect 321 221 325 224
rect 118 170 127 175
rect 150 174 154 181
rect 199 174 203 184
rect 150 169 191 174
rect 199 169 210 174
rect 313 195 317 201
rect 305 194 332 195
rect 305 190 306 194
rect 310 190 327 194
rect 331 190 332 194
rect 305 189 332 190
rect 150 166 154 169
rect 199 166 203 169
rect 135 162 172 166
rect 135 156 139 162
rect 168 156 172 162
rect 270 164 274 170
rect 262 163 289 164
rect 262 159 263 163
rect 267 159 284 163
rect 288 159 289 163
rect 262 158 289 159
rect 191 140 195 146
rect 183 139 210 140
rect 127 130 131 136
rect 160 130 164 136
rect 183 135 184 139
rect 188 135 205 139
rect 209 135 210 139
rect 183 134 210 135
rect 119 129 146 130
rect 119 125 120 129
rect 124 125 141 129
rect 145 125 146 129
rect 119 124 146 125
rect 152 129 179 130
rect 152 125 153 129
rect 157 125 174 129
rect 178 125 179 129
rect 152 124 179 125
<< labels >>
rlabel metal1 -61 254 -61 254 7 vdd
rlabel metal1 -157 254 -157 254 3 gnd
rlabel metal1 -61 305 -61 305 7 vdd
rlabel metal1 -157 305 -157 305 3 gnd
rlabel metal1 -9 247 -9 247 1 gnd
rlabel metal1 -9 343 -9 343 5 vdd
rlabel metal1 318 192 318 192 1 gnd
rlabel metal1 318 288 318 288 5 vdd
rlabel metal1 275 161 275 161 1 gnd
rlabel metal1 283 358 283 358 5 vdd
rlabel metal1 256 358 256 358 5 vdd
rlabel metal1 196 137 196 137 1 gnd
rlabel metal1 196 233 196 233 5 vdd
rlabel metal1 165 127 165 127 1 gnd
rlabel metal1 132 127 132 127 1 gnd
rlabel metal1 147 370 147 370 5 vdd
rlabel metal1 82 231 82 231 1 gnd
rlabel metal1 82 327 82 327 5 vdd
<< end >>
